package sound_pkg;

localparam int NUM_SOUNDS = 2;

localparam int Sound_Start_Length [NUM_SOUNDS][2] =
  '{'{0,    2688},
    '{2688, 30390}};

localparam int TOTOAL_LEN = Sound_Start_Length[0][1] + Sound_Start_Length[1][1];

localparam logic [11:0] Sound [TOTOAL_LEN] = {
  // ball bouncing:
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h002,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'hfff,
12'h000,
12'h002,
12'h003,
12'h000,
12'hffe,
12'h000,
12'h001,
12'h000,
12'hfff,
12'h000,
12'h003,
12'h000,
12'hfff,
12'h000,
12'h002,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'hffe,
12'h000,
12'hffd,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'hffb,
12'h000,
12'h000,
12'hffb,
12'h000,
12'h003,
12'h002,
12'h002,
12'hffc,
12'h001,
12'hfff,
12'h000,
12'hffe,
12'hffc,
12'hffe,
12'h000,
12'h002,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'hffe,
12'h000,
12'hffd,
12'hffe,
12'hffd,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'hffd,
12'hffb,
12'h000,
12'h003,
12'h001,
12'hfff,
12'h001,
12'h000,
12'h000,
12'hff9,
12'hffb,
12'h002,
12'hffc,
12'hffc,
12'h000,
12'h000,
12'h006,
12'hff9,
12'hffb,
12'hfff,
12'hff9,
12'hffe,
12'hffc,
12'h001,
12'h002,
12'h000,
12'hfff,
12'hffd,
12'h000,
12'h001,
12'hfff,
12'hfff,
12'h000,
12'h005,
12'h003,
12'h005,
12'h009,
12'hfff,
12'h006,
12'h005,
12'h004,
12'hffd,
12'h004,
12'h00d,
12'h002,
12'h000,
12'h001,
12'h000,
12'hff9,
12'hfff,
12'h002,
12'h004,
12'hffc,
12'hffc,
12'h009,
12'h001,
12'hffc,
12'hfff,
12'hffe,
12'h012,
12'hff6,
12'hff9,
12'h019,
12'h009,
12'h005,
12'h003,
12'h001,
12'h006,
12'hff4,
12'hff5,
12'h003,
12'hffd,
12'h004,
12'h005,
12'h006,
12'h005,
12'h019,
12'h015,
12'h00c,
12'h000,
12'hff9,
12'h001,
12'h00b,
12'h009,
12'h004,
12'h00d,
12'h00e,
12'h000,
12'hfff,
12'h00e,
12'h023,
12'h01a,
12'h011,
12'h031,
12'h03e,
12'h060,
12'h046,
12'h04e,
12'h0a9,
12'h0a8,
12'h051,
12'h079,
12'h0b0,
12'h111,
12'h0fd,
12'h12b,
12'h1c4,
12'h253,
12'h1ae,
12'h0d3,
12'h15f,
12'h0cd,
12'h0af,
12'h072,
12'hf1e,
12'hf77,
12'hf88,
12'hf11,
12'hf3d,
12'he20,
12'he7a,
12'he0e,
12'hdcf,
12'hdfc,
12'heac,
12'hedf,
12'hde7,
12'he5a,
12'hec4,
12'hec1,
12'hd9f,
12'hd86,
12'hd63,
12'hd92,
12'hcac,
12'hce5,
12'he1e,
12'he56,
12'hdb3,
12'hdbf,
12'hebe,
12'he2e,
12'he92,
12'hebd,
12'hf46,
12'hfc9,
12'hfc0,
12'h03d,
12'h090,
12'h0d0,
12'h10f,
12'h144,
12'h1a2,
12'h1c1,
12'h20b,
12'h2bb,
12'h33b,
12'h3c7,
12'h3b5,
12'h3e8,
12'h3ff,
12'h3a1,
12'h3ac,
12'h376,
12'h31e,
12'h28b,
12'h1e6,
12'h11e,
12'h050,
12'hfae,
12'hf16,
12'he6a,
12'he14,
12'hdf2,
12'hdc3,
12'hdad,
12'hdba,
12'hdc9,
12'hdf9,
12'he3f,
12'he5e,
12'heb3,
12'hf1a,
12'hfb0,
12'h019,
12'h07a,
12'h11c,
12'h1b3,
12'h227,
12'h2b6,
12'h2ff,
12'h306,
12'h31b,
12'h320,
12'h30c,
12'h307,
12'h2e5,
12'h249,
12'h1b0,
12'h104,
12'h028,
12'hf8e,
12'hf05,
12'he7b,
12'he26,
12'hdff,
12'hde6,
12'hdde,
12'hde5,
12'hdf1,
12'hdf4,
12'he16,
12'he7a,
12'hec1,
12'hf32,
12'hfa7,
12'h00b,
12'h084,
12'h100,
12'h17b,
12'h1cd,
12'h243,
12'h285,
12'h2a0,
12'h2b0,
12'h2b2,
12'h2c6,
12'h27d,
12'h235,
12'h1ba,
12'h114,
12'h077,
12'hfe6,
12'hf79,
12'hef6,
12'he96,
12'he5f,
12'he44,
12'he18,
12'he04,
12'he16,
12'he14,
12'he20,
12'he41,
12'he8d,
12'hee2,
12'hf23,
12'hf77,
12'hfd2,
12'h03d,
12'h0a0,
12'h101,
12'h161,
12'h1c1,
12'h1f0,
12'h20f,
12'h22c,
12'h236,
12'h22b,
12'h1f7,
12'h1aa,
12'h131,
12'h0ad,
12'h028,
12'hf9c,
12'hf14,
12'heb1,
12'he49,
12'he0f,
12'hde8,
12'hdd1,
12'hdc0,
12'hdba,
12'hdd2,
12'hde2,
12'he0c,
12'he48,
12'heac,
12'hefa,
12'hf57,
12'hfbd,
12'h020,
12'h089,
12'h0e4,
12'h12e,
12'h16b,
12'h19f,
12'h1bf,
12'h1d2,
12'h1d6,
12'h1d0,
12'h198,
12'h14d,
12'h0ee,
12'h07d,
12'h002,
12'hf82,
12'hf0e,
12'head,
12'he5f,
12'he29,
12'he09,
12'hdf5,
12'hdeb,
12'hde6,
12'hdf9,
12'he1b,
12'he43,
12'he80,
12'hed3,
12'hf24,
12'hf74,
12'hfcd,
12'h02b,
12'h07f,
12'h0c3,
12'h0fd,
12'h137,
12'h166,
12'h18a,
12'h1a2,
12'h1a7,
12'h19d,
12'h174,
12'h136,
12'h0e4,
12'h07f,
12'h015,
12'hfa7,
12'hf3c,
12'hee1,
12'he9f,
12'he6d,
12'he42,
12'he1f,
12'he0c,
12'he0d,
12'he1e,
12'he3b,
12'he68,
12'hea6,
12'heed,
12'hf37,
12'hf85,
12'hfdd,
12'h039,
12'h090,
12'h0dc,
12'h11f,
12'h15a,
12'h189,
12'h1a5,
12'h1ac,
12'h19c,
12'h17f,
12'h14e,
12'h108,
12'h0b3,
12'h058,
12'h000,
12'hfa3,
12'hf4a,
12'hefc,
12'hebf,
12'he8c,
12'he5c,
12'he3b,
12'he2c,
12'he2e,
12'he40,
12'he5e,
12'he8b,
12'hec6,
12'hf0c,
12'hf53,
12'hf9d,
12'hff2,
12'h049,
12'h09e,
12'h0ed,
12'h138,
12'h17a,
12'h1af,
12'h1ce,
12'h1d5,
12'h1c9,
12'h1ab,
12'h179,
12'h12d,
12'h0d7,
12'h07e,
12'h021,
12'hfc9,
12'hf74,
12'hf2f,
12'hef4,
12'hec0,
12'he9b,
12'he81,
12'he7d,
12'he88,
12'hea2,
12'hec7,
12'hef2,
12'hf2b,
12'hf68,
12'hfa8,
12'hfed,
12'h039,
12'h088,
12'h0d5,
12'h11b,
12'h156,
12'h186,
12'h1aa,
12'h1b9,
12'h1b6,
12'h1a1,
12'h177,
12'h13c,
12'h0f5,
12'h0a4,
12'h054,
12'hffc,
12'hfa3,
12'hf5b,
12'hf1f,
12'hef1,
12'hecb,
12'heaf,
12'hea1,
12'hea4,
12'heb7,
12'hed1,
12'hef9,
12'hf2b,
12'hf5d,
12'hf97,
12'hfd4,
12'h016,
12'h05c,
12'h09c,
12'h0e2,
12'h120,
12'h153,
12'h17e,
12'h19e,
12'h1ac,
12'h1a9,
12'h196,
12'h173,
12'h145,
12'h104,
12'h0be,
12'h071,
12'h021,
12'hfd2,
12'hf8f,
12'hf56,
12'hf21,
12'hefa,
12'hedd,
12'hed0,
12'hed2,
12'hede,
12'hef4,
12'hf19,
12'hf44,
12'hf75,
12'hfab,
12'hfe5,
12'h020,
12'h05c,
12'h099,
12'h0d2,
12'h106,
12'h133,
12'h153,
12'h16c,
12'h178,
12'h16f,
12'h156,
12'h12e,
12'h0f7,
12'h0bb,
12'h07a,
12'h037,
12'hff1,
12'hfab,
12'hf6e,
12'hf3b,
12'hf13,
12'hef7,
12'hee2,
12'hed8,
12'hedc,
12'heed,
12'hf08,
12'hf2c,
12'hf57,
12'hf8b,
12'hfc3,
12'hffb,
12'h032,
12'h06c,
12'h0a6,
12'h0dc,
12'h114,
12'h143,
12'h16a,
12'h180,
12'h187,
12'h180,
12'h165,
12'h13e,
12'h10a,
12'h0d2,
12'h093,
12'h052,
12'h010,
12'hfd4,
12'hf9a,
12'hf67,
12'hf41,
12'hf1f,
12'hf08,
12'hefc,
12'heff,
12'hf0d,
12'hf26,
12'hf43,
12'hf65,
12'hf90,
12'hfb8,
12'hfe1,
12'h00f,
12'h040,
12'h073,
12'h0a6,
12'h0d1,
12'h0fc,
12'h11c,
12'h12d,
12'h130,
12'h125,
12'h10f,
12'h0ed,
12'h0c8,
12'h09a,
12'h068,
12'h02d,
12'hff1,
12'hfb7,
12'hf7f,
12'hf4f,
12'hf29,
12'hf0f,
12'hf00,
12'hefd,
12'hf03,
12'hf10,
12'hf25,
12'hf3e,
12'hf59,
12'hf7c,
12'hfa5,
12'hfd2,
12'h004,
12'h03a,
12'h071,
12'h0a3,
12'h0d1,
12'h0f6,
12'h10f,
12'h11b,
12'h119,
12'h10e,
12'h0fb,
12'h0dd,
12'h0b9,
12'h08d,
12'h05e,
12'h029,
12'hff0,
12'hfb9,
12'hf87,
12'hf5c,
12'hf3b,
12'hf23,
12'hf16,
12'hf13,
12'hf12,
12'hf19,
12'hf27,
12'hf3f,
12'hf5a,
12'hf7b,
12'hfa3,
12'hfce,
12'hffa,
12'h027,
12'h054,
12'h07c,
12'h0a0,
12'h0be,
12'h0d6,
12'h0e1,
12'h0e3,
12'h0dc,
12'h0ca,
12'h0ac,
12'h084,
12'h05a,
12'h02e,
12'hfff,
12'hfce,
12'hf9f,
12'hf72,
12'hf4c,
12'hf30,
12'hf1b,
12'hf11,
12'hf0f,
12'hf15,
12'hf22,
12'hf38,
12'hf53,
12'hf73,
12'hf99,
12'hfbd,
12'hfe6,
12'h012,
12'h03e,
12'h065,
12'h088,
12'h0a5,
12'h0bd,
12'h0d1,
12'h0d9,
12'h0d8,
12'h0cd,
12'h0b4,
12'h094,
12'h070,
12'h047,
12'h01b,
12'hfeb,
12'hfbb,
12'hf8b,
12'hf62,
12'hf41,
12'hf28,
12'hf19,
12'hf10,
12'hf11,
12'hf1a,
12'hf28,
12'hf3d,
12'hf57,
12'hf72,
12'hf95,
12'hfbb,
12'hfe4,
12'h012,
12'h03d,
12'h066,
12'h089,
12'h0a5,
12'h0bd,
12'h0cc,
12'h0d1,
12'h0cd,
12'h0bf,
12'h0ab,
12'h08f,
12'h06d,
12'h044,
12'h017,
12'hfea,
12'hfb9,
12'hf8d,
12'hf64,
12'hf46,
12'hf2f,
12'hf20,
12'hf17,
12'hf16,
12'hf1c,
12'hf29,
12'hf3f,
12'hf58,
12'hf78,
12'hf9c,
12'hfc4,
12'hfed,
12'h017,
12'h03e,
12'h061,
12'h07e,
12'h097,
12'h0ab,
12'h0bb,
12'h0c2,
12'h0c2,
12'h0b9,
12'h0a7,
12'h08f,
12'h070,
12'h04e,
12'h02a,
12'h004,
12'hfdb,
12'hfb6,
12'hf94,
12'hf77,
12'hf5f,
12'hf4c,
12'hf3f,
12'hf3b,
12'hf3c,
12'hf46,
12'hf5a,
12'hf72,
12'hf8d,
12'hfaa,
12'hfcd,
12'hff2,
12'h018,
12'h03b,
12'h05b,
12'h077,
12'h08d,
12'h0a1,
12'h0ac,
12'h0ad,
12'h0a8,
12'h09e,
12'h08d,
12'h075,
12'h058,
12'h037,
12'h017,
12'hff2,
12'hfcc,
12'hfaa,
12'hf8b,
12'hf71,
12'hf5d,
12'hf4d,
12'hf47,
12'hf49,
12'hf51,
12'hf5b,
12'hf6b,
12'hf82,
12'hf9a,
12'hfb7,
12'hfd8,
12'hffd,
12'h01c,
12'h03d,
12'h05e,
12'h077,
12'h08d,
12'h09d,
12'h0a7,
12'h0ad,
12'h0aa,
12'h0a2,
12'h093,
12'h081,
12'h068,
12'h049,
12'h028,
12'h004,
12'hfe2,
12'hfc1,
12'hfa1,
12'hf84,
12'hf6e,
12'hf5d,
12'hf52,
12'hf50,
12'hf58,
12'hf62,
12'hf72,
12'hf86,
12'hf9d,
12'hfb8,
12'hfd8,
12'hff9,
12'h017,
12'h037,
12'h058,
12'h074,
12'h08c,
12'h09c,
12'h0a6,
12'h0a8,
12'h0a4,
12'h09b,
12'h08b,
12'h076,
12'h05d,
12'h040,
12'h021,
12'h000,
12'hfe1,
12'hfc4,
12'hfa7,
12'hf8f,
12'hf7d,
12'hf6d,
12'hf64,
12'hf62,
12'hf67,
12'hf73,
12'hf81,
12'hf95,
12'hfad,
12'hfc7,
12'hfe4,
12'h002,
12'h023,
12'h041,
12'h05e,
12'h076,
12'h08b,
12'h099,
12'h0a1,
12'h0a4,
12'h0a0,
12'h095,
12'h085,
12'h06f,
12'h057,
12'h03b,
12'h01c,
12'hffd,
12'hfdc,
12'hfbe,
12'hfa1,
12'hf8b,
12'hf79,
12'hf6c,
12'hf66,
12'hf66,
12'hf6d,
12'hf78,
12'hf87,
12'hf9a,
12'hfb1,
12'hfcc,
12'hfe8,
12'h006,
12'h023,
12'h040,
12'h05a,
12'h070,
12'h083,
12'h090,
12'h098,
12'h098,
12'h094,
12'h08b,
12'h07c,
12'h069,
12'h052,
12'h039,
12'h01c,
12'h000,
12'hfe3,
12'hfc8,
12'hfaf,
12'hf99,
12'hf88,
12'hf7c,
12'hf77,
12'hf76,
12'hf7b,
12'hf85,
12'hf93,
12'hfa4,
12'hfb8,
12'hfcf,
12'hfe8,
12'h001,
12'h01d,
12'h037,
12'h050,
12'h065,
12'h077,
12'h085,
12'h08a,
12'h08b,
12'h086,
12'h07c,
12'h06e,
12'h05c,
12'h046,
12'h02d,
12'h013,
12'hff8,
12'hfde,
12'hfc4,
12'hfad,
12'hf9a,
12'hf8b,
12'hf83,
12'hf7e,
12'hf80,
12'hf85,
12'hf8f,
12'hf9e,
12'hfae,
12'hfc2,
12'hfd9,
12'hff1,
12'h00b,
12'h024,
12'h03b,
12'h051,
12'h064,
12'h072,
12'h07e,
12'h084,
12'h084,
12'h07f,
12'h075,
12'h069,
12'h058,
12'h044,
12'h02e,
12'h016,
12'hfff,
12'hfe7,
12'hfd0,
12'hfbd,
12'hfac,
12'hf9d,
12'hf93,
12'hf8e,
12'hf8d,
12'hf92,
12'hf9b,
12'hfa8,
12'hfb7,
12'hfc9,
12'hfdf,
12'hff5,
12'h00c,
12'h024,
12'h03a,
12'h04f,
12'h05f,
12'h06e,
12'h077,
12'h07c,
12'h07a,
12'h075,
12'h06c,
12'h05f,
12'h04e,
12'h03b,
12'h026,
12'h00f,
12'hffa,
12'hfe4,
12'hfd0,
12'hfbe,
12'hfae,
12'hfa1,
12'hf99,
12'hf96,
12'hf96,
12'hf99,
12'hfa2,
12'hfad,
12'hfbb,
12'hfcb,
12'hfdc,
12'hff1,
12'h004,
12'h019,
12'h02b,
12'h03c,
12'h04c,
12'h058,
12'h060,
12'h065,
12'h066,
12'h062,
12'h05b,
12'h04f,
12'h040,
12'h032,
12'h021,
12'h00d,
12'hffb,
12'hfe8,
12'hfd7,
12'hfc6,
12'hfb8,
12'hfae,
12'hfa7,
12'hfa3,
12'hfa3,
12'hfa8,
12'hfae,
12'hfb9,
12'hfc6,
12'hfd5,
12'hfe8,
12'hffb,
12'h00f,
12'h021,
12'h033,
12'h044,
12'h052,
12'h05c,
12'h063,
12'h066,
12'h065,
12'h060,
12'h059,
12'h04e,
12'h03f,
12'h02f,
12'h01d,
12'h008,
12'hff4,
12'hfe2,
12'hfd1,
12'hfc2,
12'hfb6,
12'hfad,
12'hfa6,
12'hfa2,
12'hfa2,
12'hfa5,
12'hfab,
12'hfb5,
12'hfc1,
12'hfd0,
12'hfe1,
12'hff4,
12'h005,
12'h017,
12'h02a,
12'h039,
12'h046,
12'h050,
12'h057,
12'h05b,
12'h05c,
12'h05a,
12'h053,
12'h049,
12'h03d,
12'h02d,
12'h01c,
12'h00a,
12'hff8,
12'hfe7,
12'hfd5,
12'hfc7,
12'hfba,
12'hfb1,
12'hfaa,
12'hfa6,
12'hfa7,
12'hfab,
12'hfb1,
12'hfbc,
12'hfc9,
12'hfd7,
12'hfe9,
12'hffc,
12'h00c,
12'h01f,
12'h02f,
12'h03e,
12'h04a,
12'h053,
12'h059,
12'h05b,
12'h05a,
12'h056,
12'h04e,
12'h043,
12'h036,
12'h026,
12'h016,
12'h006,
12'hff5,
12'hfe4,
12'hfd4,
12'hfc7,
12'hfbc,
12'hfb3,
12'hfae,
12'hfab,
12'hfac,
12'hfb0,
12'hfb5,
12'hfbf,
12'hfcb,
12'hfd9,
12'hfe8,
12'hff9,
12'h009,
12'h01a,
12'h02a,
12'h038,
12'h042,
12'h04a,
12'h050,
12'h053,
12'h054,
12'h051,
12'h04b,
12'h041,
12'h035,
12'h026,
12'h016,
12'h005,
12'hff5,
12'hfe5,
12'hfd6,
12'hfc9,
12'hfbf,
12'hfb6,
12'hfb1,
12'hfaf,
12'hfb0,
12'hfb4,
12'hfba,
12'hfc4,
12'hfd0,
12'hfde,
12'hfed,
12'hffd,
12'h00b,
12'h019,
12'h027,
12'h033,
12'h03c,
12'h044,
12'h048,
12'h04a,
12'h04a,
12'h046,
12'h040,
12'h036,
12'h02a,
12'h01d,
12'h00f,
12'h000,
12'hff2,
12'hfe4,
12'hfd8,
12'hfcd,
12'hfc3,
12'hfbc,
12'hfb8,
12'hfb7,
12'hfb8,
12'hfbb,
12'hfc2,
12'hfcb,
12'hfd6,
12'hfe2,
12'hff0,
12'hffe,
12'h00b,
12'h019,
12'h025,
12'h030,
12'h03a,
12'h041,
12'h047,
12'h04a,
12'h04a,
12'h046,
12'h03f,
12'h037,
12'h02c,
12'h020,
12'h012,
12'h004,
12'hff7,
12'hfe9,
12'hfdd,
12'hfd2,
12'hfc8,
12'hfc1,
12'hfbd,
12'hfbb,
12'hfbc,
12'hfbf,
12'hfc5,
12'hfcd,
12'hfd7,
12'hfe2,
12'hfee,
12'hffa,
12'h005,
12'h011,
12'h01c,
12'h026,
12'h02e,
12'h035,
12'h038,
12'h039,
12'h038,
12'h035,
12'h02f,
12'h028,
12'h01e,
12'h014,
12'h009,
12'hffe,
12'hff3,
12'hfe8,
12'hfde,
12'hfd5,
12'hfce,
12'hfc9,
12'hfc7,
12'hfc6,
12'hfc9,
12'hfcd,
12'hfd3,
12'hfdb,
12'hfe4,
12'hfef,
12'hffb,
12'h006,
12'h011,
12'h01c,
12'h027,
12'h030,
12'h037,
12'h03d,
12'h03f,
12'h03f,
12'h03c,
12'h038,
12'h031,
12'h028,
12'h01e,
12'h012,
12'h006,
12'hffb,
12'hff0,
12'hfe5,
12'hfda,
12'hfd2,
12'hfcb,
12'hfc6,
12'hfc4,
12'hfc3,
12'hfc5,
12'hfca,
12'hfd0,
12'hfd7,
12'hfe0,
12'hfeb,
12'hff5,
12'h000,
12'h009,
12'h013,
12'h01c,
12'h025,
12'h02b,
12'h030,
12'h033,
12'h035,
12'h034,
12'h032,
12'h02d,
12'h026,
12'h01e,
12'h014,
12'h00b,
12'h001,
12'hff7,
12'hfed,
12'hfe4,
12'hfdc,
12'hfd5,
12'hfd1,
12'hfcd,
12'hfcb,
12'hfcb,
12'hfce,
12'hfd3,
12'hfda,
12'hfe1,
12'hfeb,
12'hff5,
12'hfff,
12'h008,
12'h012,
12'h01b,
12'h023,
12'h02a,
12'h02f,
12'h033,
12'h034,
12'h033,
12'h030,
12'h02b,
12'h024,
12'h01d,
12'h014,
12'h00a,
12'h000,
12'hff7,
12'hfee,
12'hfe6,
12'hfdf,
12'hfd8,
12'hfd4,
12'hfd2,
12'hfd1,
12'hfd2,
12'hfd5,
12'hfd9,
12'hfdf,
12'hfe6,
12'hff0,
12'hff9,
12'h000,
12'h008,
12'h011,
12'h01a,
12'h021,
12'h026,
12'h02a,
12'h02d,
12'h02e,
12'h02d,
12'h02b,
12'h026,
12'h020,
12'h018,
12'h010,
12'h007,
12'hffe,
12'hff5,
12'hfeb,
12'hfe3,
12'hfdd,
12'hfd6,
12'hfd2,
12'hfd0,
12'hfcf,
12'hfcf,
12'hfd2,
12'hfd8,
12'hfdf,
12'hfe6,
12'hfef,
12'hff9,
12'h002,
12'h00c,
12'h015,
12'h01d,
12'h024,
12'h029,
12'h02d,
12'h030,
12'h030,
12'h02e,
12'h02b,
12'h026,
12'h01f,
12'h018,
12'h00f,
12'h007,
12'hffe,
12'hff5,
12'hfed,
12'hfe5,
12'hfde,
12'hfd9,
12'hfd6,
12'hfd4,
12'hfd3,
12'hfd4,
12'hfd7,
12'hfdb,
12'hfe1,
12'hfe8,
12'hff0,
12'hff8,
12'h000,
12'h007,
12'h010,
12'h017,
12'h01e,
12'h023,
12'h026,
12'h028,
12'h02a,
12'h029,
12'h027,
12'h022,
12'h01d,
12'h017,
12'h010,
12'h008,
12'h000,
12'hff9,
12'hff1,
12'hfea,
12'hfe4,
12'hfdf,
12'hfdc,
12'hfda,
12'hfd9,
12'hfda,
12'hfdd,
12'hfe1,
12'hfe7,
12'hfed,
12'hff4,
12'hffb,
12'h002,
12'h00a,
12'h011,
12'h018,
12'h01d,
12'h021,
12'h024,
12'h025,
12'h025,
12'h023,
12'h020,
12'h01c,
12'h017,
12'h011,
12'h00a,
12'h003,
12'hffd,
12'hff6,
12'hfef,
12'hfe8,
12'hfe4,
12'hfe0,
12'hfdd,
12'hfdc,
12'hfdc,
12'hfdd,
12'hfe0,
12'hfe3,
12'hfe8,
12'hfed,
12'hff4,
12'hffb,
12'h001,
12'h008,
12'h00f,
12'h015,
12'h01b,
12'h01f,
12'h023,
12'h024,
12'h025,
12'h023,
12'h021,
12'h01d,
12'h018,
12'h013,
12'h00c,
12'h005,
12'hfff,
12'hff8,
12'hff1,
12'hfeb,
12'hfe7,
12'hfe2,
12'hfdf,
12'hfde,
12'hfde,
12'hfdf,
12'hfe2,
12'hfe5,
12'hfe9,
12'hfef,
12'hff5,
12'hffb,
12'h001,
12'h008,
12'h00e,
12'h013,
12'h018,
12'h01c,
12'h01e,
12'h01f,
12'h01f,
12'h01e,
12'h01b,
12'h018,
12'h014,
12'h00f,
12'h009,
12'h003,
12'hffe,
12'hff8,
12'hff2,
12'hfec,
12'hfe8,
12'hfe5,
12'hfe2,
12'hfe1,
12'hfe1,
12'hfe2,
12'hfe4,
12'hfe8,
12'hfec,
12'hff1,
12'hff7,
12'hffc,
12'h001,
12'h007,
12'h00d,
12'h013,
12'h018,
12'h01c,
12'h01e,
12'h01f,
12'h01f,
12'h01e,
12'h01b,
12'h018,
12'h014,
12'h00e,
12'h008,
12'h003,
12'hffe,
12'hff7,
12'hff1,
12'hfec,
12'hfe8,
12'hfe5,
12'hfe2,
12'hfe1,
12'hfe2,
12'hfe3,
12'hfe5,
12'hfe8,
12'hfed,
12'hff1,
12'hff6,
12'hffc,
12'h000,
12'h006,
12'h00b,
12'h010,
12'h015,
12'h018,
12'h01a,
12'h01c,
12'h01d,
12'h01c,
12'h01a,
12'h018,
12'h014,
12'h010,
12'h00b,
12'h005,
12'h000,
12'hffb,
12'hff5,
12'hff0,
12'hfeb,
12'hfe8,
12'hfe6,
12'hfe4,
12'hfe4,
12'hfe4,
12'hfe6,
12'hfe9,
12'hfed,
12'hff1,
12'hff6,
12'hffc,
12'h000,
12'h006,
12'h00b,
12'h010,
12'h014,
12'h018,
12'h01b,
12'h01c,
12'h01c,
12'h01c,
12'h01a,
12'h018,
12'h014,
12'h010,
12'h00b,
12'h006,
12'h000,
12'hffc,
12'hff6,
12'hff1,
12'hfed,
12'hfea,
12'hfe7,
12'hfe6,
12'hfe5,
12'hfe6,
12'hfe7,
12'hfea,
12'hfed,
12'hff1,
12'hff6,
12'hffa,
12'h000,
12'h004,
12'h009,
12'h00d,
12'h011,
12'h015,
12'h017,
12'h018,
12'h019,
12'h019,
12'h017,
12'h014,
12'h011,
12'h00d,
12'h008,
12'h004,
12'h000,
12'hffb,
12'hff6,
12'hff2,
12'hfee,
12'hfeb,
12'hfe8,
12'hfe7,
12'hfe7,
12'hfe8,
12'hfea,
12'hfed,
12'hff1,
12'hff5,
12'hff9,
12'hffe,
12'h002,
12'h007,
12'h00b,
12'h00f,
12'h012,
12'h015,
12'h017,
12'h018,
12'h017,
12'h016,
12'h014,
12'h011,
12'h00e,
12'h00a,
12'h006,
12'h002,
12'hffe,
12'hffa,
12'hff6,
12'hff2,
12'hfee,
12'hfec,
12'hfea,
12'hfe8,
12'hfe8,
12'hfe9,
12'hfeb,
12'hfee,
12'hff1,
12'hff5,
12'hff9,
12'hffe,
12'h002,
12'h006,
12'h00a,
12'h00e,
12'h011,
12'h013,
12'h016,
12'h017,
12'h017,
12'h016,
12'h015,
12'h013,
12'h010,
12'h00c,
12'h008,
12'h004,
12'h000,
12'hffc,
12'hff8,
12'hff4,
12'hff1,
12'hfee,
12'hfec,
12'hfeb,
12'hfeb,
12'hfeb,
12'hfed,
12'hfef,
12'hff2,
12'hff6,
12'hff9,
12'hffe,
12'h001,
12'h005,
12'h009,
12'h00c,
12'h00f,
12'h012,
12'h014,
12'h015,
12'h015,
12'h014,
12'h012,
12'h011,
12'h00e,
12'h00b,
12'h007,
12'h003,
12'h000,
12'hffc,
12'hff9,
12'hff5,
12'hff2,
12'hfef,
12'hfee,
12'hfed,
12'hfec,
12'hfed,
12'hfee,
12'hff0,
12'hff3,
12'hff6,
12'hffa,
12'hffe,
12'h000,
12'h004,
12'h008,
12'h00a,
12'h00d,
12'h010,
12'h011,
12'h012,
12'h012,
12'h011,
12'h010,
12'h00e,
12'h00b,
12'h008,
12'h005,
12'h002,
12'hfff,
12'hffc,
12'hff8,
12'hff5,
12'hff3,
12'hff1,
12'hfef,
12'hfef,
12'hfef,
12'hff0,
12'hff1,
12'hff3,
12'hff6,
12'hff9,
12'hffc,
12'hfff,
12'h002,
12'h005,
12'h009,
12'h00b,
12'h00d,
12'h00f,
12'h011,
12'h012,
12'h012,
12'h012,
12'h010,
12'h00f,
12'h00c,
12'h00a,
12'h006,
12'h003,
12'h000,
12'hffd,
12'hffa,
12'hff7,
12'hff4,
12'hff2,
12'hff0,
12'hfef,
12'hfee,
12'hfef,
12'hff0,
12'hff1,
12'hff4,
12'hff6,
12'hff9,
12'hffc,
12'h000,
12'h002,
12'h005,
12'h008,
12'h00a,
12'h00c,
12'h00e,
12'h00f,
12'h00f,
12'h00f,
12'h00e,
12'h00d,
12'h00b,
12'h009,
12'h006,
12'h003,
12'h000,
12'hffe,
12'hffb,
12'hff8,
12'hff6,
12'hff4,
12'hff3,
12'hff2,
12'hff2,
12'hff2,
12'hff3,
12'hff5,
12'hff6,
12'hff9,
12'hffb,
12'hffe,
12'h000,
12'h003,
12'h005,
12'h008,
12'h00a,
12'h00c,
12'h00d,
12'h00e,
12'h00f,
12'h00e,
12'h00e,
12'h00d,
12'h00b,
12'h009,
12'h006,
12'h004,
12'h001,
12'hfff,
12'hffc,
12'hff9,
12'hff7,
12'hff5,
12'hff3,
12'hff2,
12'hff2,
12'hff2,
12'hff3,
12'hff4,
12'hff6,
12'hff8,
12'hffb,
12'hffd,
12'h000,
12'h001,
12'h004,
12'h006,
12'h009,
12'h00a,
12'h00b,
12'h00c,
12'h00c,
12'h00c,
12'h00c,
12'h00b,
12'h009,
12'h007,
12'h005,
12'h003,
12'h000,
12'hfff,
12'hffc,
12'hffa,
12'hff8,
12'hff6,
12'hff5,
12'hff4,
12'hff4,
12'hff4,
12'hff5,
12'hff6,
12'hff7,
12'hff9,
12'hffb,
12'hffe,
12'h000,
12'h002,
12'h004,
12'h006,
12'h007,
12'h009,
12'h00b,
12'h00b,
12'h00c,
12'h00c,
12'h00b,
12'h00a,
12'h009,
12'h007,
12'h004,
12'h002,
12'h000,
12'hffe,
12'hffc,
12'hffa,
12'hff8,
12'hff7,
12'hff6,
12'hff5,
12'hff5,
12'hff5,
12'hff6,
12'hff8,
12'hff9,
12'hffb,
12'hffe,
12'h000,
12'h001,
12'h003,
12'h005,
12'h007,
12'h009,
12'h00a,
12'h00a,
12'h00a,
12'h00b,
12'h00b,
12'h00a,
12'h009,
12'h008,
12'h006,
12'h004,
12'h002,
12'h000,
12'hfff,
12'hffd,
12'hffb,
12'hffa,
12'hff8,
12'hff7,
12'hff6,
12'hff6,
12'hff6,
12'hff7,
12'hff7,
12'hff9,
12'hffa,
12'hffc,
12'hffe,
12'h000,
12'h001,
12'h003,
12'h004,
12'h006,
12'h007,
12'h008,
12'h009,
12'h009,
12'h009,
12'h008,
12'h007,
12'h006,
12'h005,
12'h003,
12'h001,
12'h000,
12'hffe,
12'hffd,
12'hffb,
12'hff9,
12'hff8,
12'hff7,
12'hff7,
12'hff7,
12'hff7,
12'hff8,
12'hff9,
12'hffa,
12'hffc,
12'hffe,
12'hfff,
12'h000,
12'h002,
12'h004,
12'h005,
12'h006,
12'h008,
12'h008,
12'h009,
12'h009,
12'h009,
12'h009,
12'h008,
12'h008,
12'h006,
12'h005,
12'h003,
12'h002,
12'h000,
12'hfff,
12'hffd,
12'hffc,
12'hffa,
12'hff8,
12'hff7,
12'hff7,
12'hff7,
12'hff7,
12'hff8,
12'hff9,
12'hffb,
12'hffc,
12'hffe,
12'hfff,
12'h000,
12'h002,
12'h004,
12'h005,
12'h006,
12'h007,
12'h008,
12'h008,
12'h008,
12'h008,
12'h007,
12'h006,
12'h005,
12'h004,
12'h003,
12'h001,
12'h000,
12'hfff,
12'hffd,
12'hffc,
12'hffb,
12'hffa,
12'hff9,
12'hff9,
12'hff9,
12'hffa,
12'hffa,
12'hffb,
12'hffc,
12'hffc,
12'hffe,
12'hfff,
12'h000,
12'h001,
12'h002,
12'h003,
12'h004,
12'h005,
12'h006,
12'h006,
12'h007,
12'h007,
12'h006,
12'h006,
12'h005,
12'h004,
12'h003,
12'h001,
12'h000,
12'h000,
12'hffe,
12'hffd,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffc,
12'hffd,
12'hffd,
12'hffe,
12'h000,
12'h000,
12'h000,
12'h001,
12'h002,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h002,
12'h002,
12'h001,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hffe,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffe,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h001,
12'h002,
12'h003,
12'h004,
12'h004,
12'h005,
12'h005,
12'h005,
12'h005,
12'h004,
12'h004,
12'h003,
12'h002,
12'h001,
12'h000,
12'h000,
12'hfff,
12'hffe,
12'hffd,
12'hffc,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffd,
12'hffe,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'h001,
12'h002,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h002,
12'h002,
12'h001,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'hffe,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffe,
12'hfff,
12'h000,
12'h000,
12'h001,
12'h002,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h002,
12'h001,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'hffe,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h002,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'hffe,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h001,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hffe,
12'hffe,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hffe,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'hfff,
12'hffe,
12'hffe,
12'hffe,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
// End Game

12'hfff,
12'hffd,
12'hffa,
12'hffa,
12'hffa,
12'hffb,
12'hffb,
12'hffb,
12'hffa,
12'hffa,
12'hffa,
12'hffa,
12'hffa,
12'hffa,
12'hffb,
12'hffb,
12'hffa,
12'hffa,
12'hffa,
12'hffa,
12'hffa,
12'hffc,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hffd,
12'hffa,
12'hff9,
12'hffa,
12'hffa,
12'hffa,
12'hffa,
12'hffa,
12'hffc,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hffc,
12'hffa,
12'hffa,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffd,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'h000,
12'h005,
12'h00b,
12'h00c,
12'h007,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hffe,
12'hffb,
12'hff9,
12'hffa,
12'hffb,
12'hffb,
12'hffa,
12'hffb,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'h000,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'h000,
12'h000,
12'hfff,
12'hffe,
12'hfff,
12'h000,
12'h001,
12'h001,
12'h001,
12'h002,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h000,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hffe,
12'hffc,
12'hff9,
12'hff8,
12'hff8,
12'hffa,
12'hffb,
12'hffc,
12'hffd,
12'hfff,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'hfff,
12'hffe,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'hfff,
12'hffe,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h001,
12'h002,
12'h000,
12'h000,
12'h000,
12'hffe,
12'hffc,
12'hffb,
12'hff9,
12'hff8,
12'hff6,
12'hff5,
12'hff6,
12'hff9,
12'hffa,
12'hffa,
12'hffc,
12'hfff,
12'h000,
12'h001,
12'h002,
12'h003,
12'h003,
12'h001,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h001,
12'h001,
12'h001,
12'h002,
12'h001,
12'h000,
12'hffd,
12'hff9,
12'hff7,
12'hff8,
12'hffa,
12'hffd,
12'h000,
12'h002,
12'h001,
12'h000,
12'h001,
12'h000,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h003,
12'h003,
12'h001,
12'h000,
12'h005,
12'h009,
12'h00b,
12'h00c,
12'h00c,
12'h006,
12'h000,
12'h000,
12'h003,
12'h005,
12'h004,
12'h002,
12'h000,
12'h000,
12'hffe,
12'hffb,
12'hff9,
12'hff7,
12'hff5,
12'hff1,
12'hff0,
12'hff1,
12'hff0,
12'hfed,
12'hfef,
12'hff2,
12'hff2,
12'hff3,
12'hff7,
12'hff9,
12'hff9,
12'hffb,
12'hffe,
12'hffe,
12'hffe,
12'h000,
12'h000,
12'hfff,
12'hfff,
12'h000,
12'h000,
12'hfff,
12'h000,
12'h001,
12'h001,
12'h000,
12'h001,
12'h002,
12'h003,
12'h004,
12'h003,
12'h002,
12'h001,
12'h002,
12'h005,
12'h006,
12'h007,
12'h006,
12'h005,
12'h007,
12'h00b,
12'h011,
12'h015,
12'h013,
12'h010,
12'h00e,
12'h00e,
12'h00d,
12'h00c,
12'h00b,
12'h006,
12'h000,
12'hffc,
12'hffd,
12'hffe,
12'hfff,
12'h000,
12'hffe,
12'hffc,
12'hffc,
12'hfff,
12'h000,
12'hfff,
12'hffe,
12'hffb,
12'hff7,
12'hff4,
12'hff3,
12'hff2,
12'hfee,
12'hfea,
12'hfe4,
12'hfe0,
12'hfdd,
12'hfdd,
12'hfdd,
12'hfde,
12'hfe1,
12'hfe3,
12'hfe6,
12'hfed,
12'hff4,
12'hffa,
12'hffd,
12'h000,
12'h000,
12'h001,
12'h005,
12'h00b,
12'h00e,
12'h00e,
12'h00e,
12'h00c,
12'h00b,
12'h00d,
12'h010,
12'h011,
12'h00e,
12'h00a,
12'h006,
12'h003,
12'h002,
12'h003,
12'h004,
12'h002,
12'h001,
12'h001,
12'h002,
12'h003,
12'h004,
12'h003,
12'h002,
12'h000,
12'hffe,
12'hffd,
12'hffe,
12'hffe,
12'hfff,
12'hfff,
12'hfff,
12'hffe,
12'hfff,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hffd,
12'hffa,
12'hff9,
12'hffa,
12'hffe,
12'h000,
12'h001,
12'h001,
12'h000,
12'hfff,
12'hffd,
12'hffa,
12'hff6,
12'hff1,
12'hfeb,
12'hfe7,
12'hfe3,
12'hfe2,
12'hfe3,
12'hfe5,
12'hfe9,
12'hfed,
12'hff1,
12'hff6,
12'hffa,
12'hffd,
12'hfff,
12'h000,
12'h001,
12'h004,
12'h00a,
12'h010,
12'h016,
12'h01b,
12'h01e,
12'h01e,
12'h01e,
12'h01d,
12'h01b,
12'h019,
12'h013,
12'h00e,
12'h008,
12'h004,
12'h001,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h001,
12'h002,
12'h001,
12'h000,
12'h000,
12'hffe,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hfff,
12'hfff,
12'hffe,
12'h000,
12'h001,
12'h002,
12'h000,
12'h000,
12'h000,
12'hffe,
12'hffe,
12'h000,
12'h002,
12'h001,
12'h000,
12'h000,
12'hfff,
12'hffe,
12'h000,
12'h000,
12'hfff,
12'hffe,
12'hffc,
12'hffa,
12'hffa,
12'hffd,
12'h000,
12'h003,
12'h006,
12'h006,
12'h005,
12'h004,
12'h004,
12'h003,
12'h003,
12'h004,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h000,
12'hfff,
12'hfff,
12'h001,
12'h002,
12'h001,
12'hfff,
12'hffc,
12'hffb,
12'hffa,
12'hffb,
12'hffc,
12'hffe,
12'hfff,
12'hfff,
12'hffd,
12'hffc,
12'hffe,
12'hfff,
12'h001,
12'h001,
12'h000,
12'hfff,
12'hffe,
12'hffe,
12'hffd,
12'hffc,
12'hffb,
12'hffe,
12'hfff,
12'hfff,
12'h000,
12'h001,
12'h001,
12'h003,
12'h006,
12'h006,
12'h004,
12'h003,
12'h002,
12'h001,
12'h002,
12'h001,
12'h001,
12'h004,
12'h001,
12'hffe,
12'hff8,
12'hff1,
12'hfea,
12'hfe3,
12'hfe2,
12'hfe4,
12'hfe6,
12'hfe4,
12'hfef,
12'hffd,
12'hffd,
12'h000,
12'h006,
12'h00b,
12'h00b,
12'h00c,
12'h00d,
12'h00e,
12'h009,
12'h002,
12'h005,
12'h000,
12'hffc,
12'hffa,
12'hffa,
12'hff7,
12'hff4,
12'hff7,
12'hff6,
12'hff6,
12'hff7,
12'hff9,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hff8,
12'hff6,
12'hff6,
12'hff7,
12'hff4,
12'hff2,
12'hff2,
12'hff2,
12'hff3,
12'hff5,
12'hff9,
12'hffe,
12'h000,
12'h000,
12'h003,
12'h006,
12'h009,
12'h009,
12'h002,
12'hffb,
12'hffb,
12'hffc,
12'hffd,
12'hffe,
12'hffb,
12'hffd,
12'hfff,
12'h000,
12'h004,
12'h008,
12'h008,
12'h002,
12'hff9,
12'hff2,
12'hfee,
12'hfe7,
12'hfe3,
12'hfe6,
12'hfec,
12'hff1,
12'hff4,
12'hff6,
12'hff6,
12'hff6,
12'hff8,
12'hffd,
12'hffc,
12'hff5,
12'hfef,
12'hfee,
12'hff2,
12'hff7,
12'hffe,
12'h002,
12'h007,
12'h00a,
12'h011,
12'h014,
12'h00e,
12'h006,
12'h000,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'h001,
12'h00a,
12'h00d,
12'h011,
12'h017,
12'h01a,
12'h014,
12'h00b,
12'h00b,
12'h016,
12'h01c,
12'h013,
12'h005,
12'h000,
12'h002,
12'hffc,
12'hff6,
12'hffe,
12'h010,
12'h01c,
12'h016,
12'h014,
12'h025,
12'h033,
12'h02e,
12'h025,
12'h031,
12'h04b,
12'h052,
12'h03f,
12'h028,
12'h01e,
12'h020,
12'h015,
12'hffb,
12'hfc6,
12'hf71,
12'hf15,
12'hecd,
12'hebd,
12'hedf,
12'hf16,
12'hf54,
12'hf91,
12'hfcf,
12'h010,
12'h04f,
12'h06c,
12'h04b,
12'hffb,
12'hf9a,
12'hf53,
12'hf2e,
12'hf20,
12'hf24,
12'hf2e,
12'hf44,
12'hf84,
12'hff2,
12'h075,
12'h0ce,
12'h0c9,
12'h07b,
12'h012,
12'hfb0,
12'hf73,
12'hf82,
12'hfd0,
12'h022,
12'h04c,
12'h044,
12'h048,
12'h07f,
12'h0c1,
12'h0f0,
12'h0fe,
12'h0ed,
12'h0c1,
12'h085,
12'h058,
12'h04a,
12'h050,
12'h055,
12'h065,
12'h08b,
12'h0b9,
12'h0ce,
12'h0d7,
12'h0f2,
12'h106,
12'h0fc,
12'h0d1,
12'h0a6,
12'h088,
12'h060,
12'h043,
12'h043,
12'h067,
12'h086,
12'h075,
12'h047,
12'h02b,
12'h02b,
12'h02a,
12'h017,
12'hff2,
12'hfda,
12'hfda,
12'hfef,
12'h023,
12'h065,
12'h08b,
12'h06a,
12'h025,
12'hffa,
12'hff3,
12'hfe7,
12'hfc5,
12'hfad,
12'hfab,
12'hfb1,
12'hfae,
12'hfb1,
12'hfb9,
12'hfae,
12'hf9c,
12'hf91,
12'hfa8,
12'hfd4,
12'hff1,
12'hff3,
12'hfe1,
12'hfd0,
12'hfb8,
12'hf92,
12'hf5d,
12'hf3a,
12'hf2f,
12'hf2b,
12'hf3e,
12'hf6f,
12'hfb1,
12'hfe1,
12'hffc,
12'h009,
12'h007,
12'hfe2,
12'hf9e,
12'hf67,
12'hf54,
12'hf67,
12'hf96,
12'hfc9,
12'hfd1,
12'hfac,
12'hf89,
12'hf7a,
12'hf7d,
12'hf92,
12'hfc3,
12'hff7,
12'hfff,
12'hfd3,
12'hfa7,
12'hf9f,
12'hfa9,
12'hfac,
12'hfb7,
12'hfd9,
12'hffa,
12'hffe,
12'hff3,
12'hfef,
12'hffa,
12'h006,
12'h005,
12'hffb,
12'hfe7,
12'hfd2,
12'hfc4,
12'hfc5,
12'hfdb,
12'hffa,
12'h00a,
12'h00a,
12'h007,
12'h00d,
12'h017,
12'h011,
12'h007,
12'h012,
12'h028,
12'h03f,
12'h050,
12'h065,
12'h087,
12'h0a2,
12'h0a5,
12'h092,
12'h06d,
12'h045,
12'h02e,
12'h023,
12'h02c,
12'h04f,
12'h086,
12'h0b5,
12'h0d0,
12'h0d8,
12'h0c8,
12'h0b2,
12'h09e,
12'h08c,
12'h084,
12'h091,
12'h0a2,
12'h0a8,
12'h0ac,
12'h0b0,
12'h0b1,
12'h0ac,
12'h0a3,
12'h0a1,
12'h0a1,
12'h090,
12'h066,
12'h03e,
12'h039,
12'h04c,
12'h063,
12'h072,
12'h07c,
12'h078,
12'h065,
12'h04a,
12'h037,
12'h045,
12'h06a,
12'h085,
12'h07e,
12'h069,
12'h066,
12'h075,
12'h073,
12'h05f,
12'h050,
12'h042,
12'h02b,
12'h00e,
12'hff6,
12'hfe9,
12'hfdf,
12'hfce,
12'hfb9,
12'hfab,
12'hfa4,
12'hf92,
12'hf70,
12'hf52,
12'hf46,
12'hf50,
12'hf6a,
12'hf93,
12'hfc4,
12'hfd3,
12'hfae,
12'hf77,
12'hf60,
12'hf73,
12'hf85,
12'hf7e,
12'hf79,
12'hf92,
12'hfaa,
12'hf8d,
12'hf45,
12'hf0c,
12'heed,
12'hec2,
12'he73,
12'he20,
12'hdf6,
12'he00,
12'he30,
12'he72,
12'hec1,
12'hf08,
12'hf1c,
12'hefe,
12'hee3,
12'hee1,
12'heea,
12'heda,
12'heab,
12'he90,
12'he94,
12'heb4,
12'hef5,
12'hf4b,
12'hfa8,
12'hfda,
12'hfad,
12'hf40,
12'hedd,
12'heb1,
12'heb2,
12'hec6,
12'heea,
12'hf0b,
12'hf1b,
12'hf32,
12'hf72,
12'h000,
12'h099,
12'h0d9,
12'h0ab,
12'h03f,
12'hff2,
12'hfde,
12'h000,
12'h05c,
12'h0f6,
12'h19f,
12'h1e2,
12'h1d4,
12'h1cb,
12'h1e8,
12'h20c,
12'h1f4,
12'h1bb,
12'h189,
12'h172,
12'h19b,
12'h1f1,
12'h24b,
12'h277,
12'h25f,
12'h225,
12'h1e6,
12'h1a6,
12'h16e,
12'h156,
12'h16b,
12'h18f,
12'h19e,
12'h19e,
12'h1a2,
12'h1b3,
12'h1c0,
12'h1c3,
12'h1c3,
12'h1a9,
12'h16f,
12'h115,
12'h0c5,
12'h0ab,
12'h0ac,
12'h094,
12'h034,
12'hfc3,
12'hf92,
12'hf9c,
12'hfd0,
12'h016,
12'h071,
12'h0b5,
12'h096,
12'h028,
12'hfaf,
12'hf68,
12'hf4a,
12'hf33,
12'hf2b,
12'hf42,
12'hf66,
12'hf6d,
12'hf54,
12'hf2f,
12'hf1a,
12'hf0c,
12'hedf,
12'heaa,
12'he95,
12'he9f,
12'heb1,
12'hec8,
12'hee9,
12'hf1f,
12'hf4e,
12'hf57,
12'hf42,
12'hf19,
12'heed,
12'hecd,
12'hecf,
12'heff,
12'hf44,
12'hf5f,
12'hf45,
12'hf12,
12'heea,
12'hee4,
12'hef0,
12'hf01,
12'hf1d,
12'hf46,
12'hf6e,
12'hf7e,
12'hf80,
12'hfa5,
12'hff3,
12'h04e,
12'h07f,
12'h076,
12'h068,
12'h06e,
12'h07d,
12'h097,
12'h0be,
12'h0cf,
12'h0b6,
12'h076,
12'h033,
12'h024,
12'h04b,
12'h085,
12'h0ad,
12'h0a1,
12'h085,
12'h088,
12'h0b1,
12'h0f3,
12'h128,
12'h133,
12'h111,
12'h0d1,
12'h08b,
12'h055,
12'h048,
12'h070,
12'h0a7,
12'h0be,
12'h0a8,
12'h078,
12'h056,
12'h055,
12'h05e,
12'h060,
12'h054,
12'h02d,
12'hffb,
12'hfcc,
12'hfa3,
12'hf87,
12'hf78,
12'hf6d,
12'hf5a,
12'hf2d,
12'hf05,
12'hf0a,
12'hf3c,
12'hf7d,
12'hfa1,
12'hf9e,
12'hf7d,
12'hf47,
12'hf0b,
12'hed2,
12'heac,
12'hea8,
12'hec0,
12'hf02,
12'hf57,
12'hfa3,
12'hfbc,
12'hf81,
12'hf1a,
12'hec6,
12'he90,
12'he4c,
12'hdfb,
12'hdc2,
12'hdd9,
12'he4a,
12'hec6,
12'hef4,
12'hedb,
12'heb7,
12'hea9,
12'he97,
12'he75,
12'he62,
12'he67,
12'he6f,
12'he7e,
12'hec5,
12'hf58,
12'hff7,
12'h036,
12'hff2,
12'hf6c,
12'hf13,
12'hf1b,
12'hf74,
12'hfe1,
12'h020,
12'h015,
12'hffb,
12'h011,
12'h05a,
12'h0b0,
12'h0e2,
12'h0ef,
12'h0d2,
12'h088,
12'h048,
12'h060,
12'h0d3,
12'h159,
12'h1b1,
12'h1dc,
12'h1ff,
12'h234,
12'h263,
12'h281,
12'h2a6,
12'h2b5,
12'h272,
12'h1f4,
12'h199,
12'h192,
12'h1c9,
12'h1f9,
12'h209,
12'h200,
12'h1ee,
12'h1eb,
12'h200,
12'h220,
12'h215,
12'h1d2,
12'h163,
12'h0dd,
12'h05e,
12'h00e,
12'h018,
12'h077,
12'h0fc,
12'h162,
12'h18c,
12'h181,
12'h13e,
12'h0d8,
12'h061,
12'hfee,
12'hf8f,
12'hf54,
12'hf48,
12'hf5c,
12'hf7f,
12'hfa5,
12'hfba,
12'hfba,
12'hfa1,
12'hf5e,
12'hf03,
12'heb3,
12'he87,
12'he7f,
12'he91,
12'heb2,
12'hecf,
12'hee8,
12'hef6,
12'hee1,
12'head,
12'he72,
12'he4c,
12'he45,
12'he64,
12'he96,
12'hec2,
12'hedd,
12'hee4,
12'hef4,
12'hf24,
12'hf51,
12'hf52,
12'hf31,
12'hf1b,
12'hf38,
12'hf70,
12'hfa0,
12'hfd1,
12'h009,
12'h026,
12'h00c,
12'hfe2,
12'hfcd,
12'hfcd,
12'hfe0,
12'h002,
12'h025,
12'h041,
12'h04b,
12'h04b,
12'h056,
12'h07a,
12'h0a8,
12'h0df,
12'h119,
12'h12f,
12'h128,
12'h11a,
12'h11d,
12'h133,
12'h13d,
12'h137,
12'h12f,
12'h130,
12'h12e,
12'h121,
12'h11b,
12'h10c,
12'h0e6,
12'h0a9,
12'h076,
12'h076,
12'h096,
12'h0bd,
12'h0df,
12'h0fd,
12'h10b,
12'h0fd,
12'h0ee,
12'h0eb,
12'h0f3,
12'h0df,
12'h0a3,
12'h07d,
12'h06f,
12'h064,
12'h058,
12'h04b,
12'h05a,
12'h066,
12'h05a,
12'h036,
12'h000,
12'hfcc,
12'hf7f,
12'hf23,
12'hed6,
12'hea0,
12'he93,
12'hea2,
12'heac,
12'hea7,
12'heaf,
12'hed9,
12'hf09,
12'hf06,
12'heb5,
12'he65,
12'he4d,
12'he48,
12'he26,
12'hdee,
12'hde7,
12'he2b,
12'he7f,
12'hea4,
12'hea7,
12'heb6,
12'hecf,
12'hec2,
12'he92,
12'he5e,
12'he3d,
12'he35,
12'he20,
12'hdfd,
12'hde6,
12'hdf2,
12'he2b,
12'he73,
12'heb0,
12'hee0,
12'hef7,
12'heee,
12'hec6,
12'heb3,
12'hedf,
12'hf30,
12'hf80,
12'hfb2,
12'hfda,
12'hffb,
12'hfff,
12'hfe4,
12'hfbe,
12'hf9e,
12'hf7a,
12'hf4b,
12'hf2e,
12'hf4d,
12'hfb0,
12'h03c,
12'h0e7,
12'h17c,
12'h199,
12'h140,
12'h0d2,
12'h0b0,
12'h0d6,
12'h0fb,
12'h0e8,
12'h0d0,
12'h10a,
12'h179,
12'h1fa,
12'h292,
12'h336,
12'h3af,
12'h3a0,
12'h319,
12'h27f,
12'h224,
12'h210,
12'h20c,
12'h207,
12'h1fe,
12'h1fc,
12'h21d,
12'h263,
12'h29b,
12'h2ad,
12'h29a,
12'h271,
12'h234,
12'h1e8,
12'h1b2,
12'h18d,
12'h15e,
12'h11c,
12'h0e2,
12'h0d1,
12'h0e8,
12'h118,
12'h13c,
12'h137,
12'h10f,
12'h0c2,
12'h062,
12'h01c,
12'hff7,
12'hfe2,
12'hfdf,
12'hfe5,
12'hfea,
12'hfdd,
12'hfb8,
12'hf86,
12'hf5e,
12'hf2f,
12'hef0,
12'hec2,
12'hea8,
12'he9e,
12'he9f,
12'hebc,
12'heef,
12'hf06,
12'hefb,
12'hedb,
12'hec7,
12'hebf,
12'hea9,
12'he8f,
12'he6c,
12'he54,
12'he53,
12'he57,
12'he59,
12'he5a,
12'he68,
12'he7c,
12'he89,
12'he96,
12'heae,
12'hee8,
12'hf3a,
12'hf70,
12'hf73,
12'hf43,
12'hef4,
12'heb3,
12'hea8,
12'heca,
12'hee8,
12'hef5,
12'hf00,
12'hf1f,
12'hf4e,
12'hf86,
12'hfc6,
12'hff9,
12'h019,
12'h02d,
12'h03f,
12'h06c,
12'h0b4,
12'h0fb,
12'h115,
12'h0ff,
12'h0e6,
12'h0df,
12'h0eb,
12'h0f7,
12'h105,
12'h114,
12'h11f,
12'h12e,
12'h137,
12'h146,
12'h15c,
12'h158,
12'h12f,
12'h0e9,
12'h0ac,
12'h0a9,
12'h0d2,
12'h102,
12'h12c,
12'h144,
12'h149,
12'h130,
12'h0ff,
12'h0ce,
12'h0a1,
12'h08b,
12'h084,
12'h07a,
12'h05e,
12'h049,
12'h044,
12'h044,
12'h041,
12'h030,
12'h002,
12'hfa4,
12'hf2d,
12'hecc,
12'heac,
12'hed3,
12'hf1a,
12'hf54,
12'hf6e,
12'hf50,
12'hf02,
12'hebe,
12'heab,
12'heba,
12'heb0,
12'he7b,
12'he34,
12'he04,
12'he02,
12'he1a,
12'he57,
12'heac,
12'hedc,
12'hec8,
12'hea0,
12'head,
12'heeb,
12'hf21,
12'hf27,
12'hf15,
12'hef9,
12'hec6,
12'he79,
12'he37,
12'he46,
12'he8e,
12'hec2,
12'heca,
12'hec8,
12'hed3,
12'heef,
12'hf21,
12'hf61,
12'hfa5,
12'hfcf,
12'hfba,
12'hf75,
12'hf25,
12'hefa,
12'hf06,
12'hf2b,
12'hf4d,
12'hf4c,
12'hf30,
12'hf27,
12'hf5e,
12'hfda,
12'h070,
12'h0d0,
12'h0c3,
12'h067,
12'hfed,
12'hf89,
12'hf72,
12'hfa4,
12'hfe7,
12'h008,
12'h011,
12'h02a,
12'h07e,
12'h104,
12'h193,
12'h1f1,
12'h205,
12'h1d0,
12'h161,
12'h0f9,
12'h0e2,
12'h140,
12'h1db,
12'h275,
12'h2cf,
12'h2eb,
12'h301,
12'h30e,
12'h303,
12'h2cc,
12'h282,
12'h246,
12'h218,
12'h213,
12'h226,
12'h24d,
12'h27b,
12'h289,
12'h265,
12'h213,
12'h1bc,
12'h17e,
12'h162,
12'h162,
12'h15a,
12'h148,
12'h136,
12'h114,
12'h0e9,
12'h0c7,
12'h0c2,
12'h0d5,
12'h0da,
12'h0c2,
12'h075,
12'h000,
12'hf90,
12'hf3a,
12'heff,
12'hec9,
12'hea8,
12'heb5,
12'hed0,
12'hee3,
12'heee,
12'hf09,
12'hf39,
12'hf65,
12'hf75,
12'hf54,
12'hf0a,
12'head,
12'he4e,
12'he12,
12'he19,
12'he6f,
12'hee2,
12'hf2b,
12'hf2f,
12'hf01,
12'hed4,
12'hec8,
12'hee3,
12'hf09,
12'hf16,
12'hf11,
12'hf02,
12'hf02,
12'hf2d,
12'hf7d,
12'hfda,
12'h013,
12'hffd,
12'hf97,
12'hf2b,
12'hefb,
12'hf1d,
12'hf7a,
12'hfdb,
12'h006,
12'hfe6,
12'hfa5,
12'hf7a,
12'hf72,
12'hf95,
12'hfd4,
12'h006,
12'h011,
12'hfdd,
12'hf92,
12'hf88,
12'hfe9,
12'h08e,
12'h108,
12'h121,
12'h0ed,
12'h09c,
12'h06c,
12'h06e,
12'h0b0,
12'h10e,
12'h133,
12'h101,
12'h099,
12'h05d,
12'h070,
12'h0a4,
12'h0c5,
12'h0b2,
12'h080,
12'h03f,
12'h009,
12'h01e,
12'h076,
12'h0d5,
12'h0f5,
12'h0ac,
12'h027,
12'hfb3,
12'hf7e,
12'hf93,
12'hfce,
12'h012,
12'h037,
12'h020,
12'hfe8,
12'hfb4,
12'hfa1,
12'hfad,
12'hfb3,
12'hf9f,
12'hf7c,
12'hf4c,
12'hf07,
12'hebe,
12'he8a,
12'he76,
12'he6b,
12'he4a,
12'he29,
12'he2c,
12'he51,
12'he87,
12'hecd,
12'hf20,
12'hf57,
12'hf4a,
12'hf05,
12'hec2,
12'he97,
12'he74,
12'he50,
12'he60,
12'hec9,
12'hf4d,
12'hf9e,
12'hfa8,
12'hf89,
12'hf61,
12'hf2c,
12'hee4,
12'he9c,
12'he76,
12'he7b,
12'heab,
12'hf05,
12'hf81,
12'h002,
12'h05a,
12'h060,
12'h013,
12'hf9b,
12'hf2f,
12'hef2,
12'hed5,
12'hed5,
12'hf0d,
12'hf8b,
12'h03c,
12'h0db,
12'h151,
12'h1ab,
12'h1c7,
12'h18f,
12'h0fe,
12'h06e,
12'h02d,
12'h008,
12'hff8,
12'h012,
12'h05d,
12'h0d4,
12'h160,
12'h1fe,
12'h282,
12'h2c3,
12'h2d5,
12'h2bf,
12'h292,
12'h244,
12'h1bd,
12'h128,
12'h0cf,
12'h0ee,
12'h17e,
12'h235,
12'h2d8,
12'h33c,
12'h35f,
12'h355,
12'h32b,
12'h2fb,
12'h2b6,
12'h258,
12'h1f1,
12'h191,
12'h145,
12'h0ff,
12'h0d4,
12'h0d2,
12'h0f1,
12'h130,
12'h172,
12'h199,
12'h194,
12'h156,
12'h0f1,
12'h079,
12'h010,
12'hfe5,
12'h003,
12'h02e,
12'h01d,
12'hfcb,
12'hf60,
12'hf1e,
12'hf01,
12'hedf,
12'heb4,
12'he82,
12'he5f,
12'he65,
12'he95,
12'hedd,
12'hef7,
12'hec5,
12'he62,
12'hdfa,
12'hdb2,
12'hd95,
12'hdab,
12'hdd9,
12'hdfa,
12'he04,
12'hdf6,
12'hde6,
12'hde3,
12'hdfe,
12'he33,
12'he68,
12'he8a,
12'he7e,
12'he4e,
12'he21,
12'he10,
12'he34,
12'he83,
12'hed1,
12'hef0,
12'hee0,
12'hec9,
12'hecb,
12'hee1,
12'hf0a,
12'hf5a,
12'hfc1,
12'h008,
12'h01a,
12'h021,
12'h03f,
12'h05f,
12'h062,
12'h047,
12'h022,
12'hffb,
12'hfe3,
12'hff1,
12'h032,
12'h097,
12'h0dc,
12'h107,
12'h142,
12'h187,
12'h1c5,
12'h1ed,
12'h215,
12'h23b,
12'h242,
12'h227,
12'h1eb,
12'h1bc,
12'h1a4,
12'h18a,
12'h17b,
12'h190,
12'h1bf,
12'h1e3,
12'h1e6,
12'h1d0,
12'h1b1,
12'h18b,
12'h16b,
12'h167,
12'h162,
12'h147,
12'h116,
12'h0e5,
12'h0c5,
12'h0ba,
12'h0d2,
12'h0e8,
12'h0f3,
12'h0eb,
12'h0b2,
12'h064,
12'h016,
12'hfee,
12'hfeb,
12'hffc,
12'h008,
12'hff8,
12'hfd0,
12'hf87,
12'hf39,
12'hefb,
12'heb9,
12'he71,
12'he10,
12'hdac,
12'hd7b,
12'hd90,
12'hddb,
12'he34,
12'he7d,
12'hea0,
12'he94,
12'he66,
12'he29,
12'hdea,
12'hdbe,
12'hdcf,
12'he05,
12'he25,
12'he27,
12'he22,
12'he39,
12'he7e,
12'hec2,
12'hed3,
12'hecc,
12'hec2,
12'he95,
12'he3a,
12'hdd9,
12'hdc2,
12'he02,
12'he68,
12'hed7,
12'hf36,
12'hf79,
12'hf9a,
12'hfa3,
12'hfa1,
12'hfae,
12'hfbe,
12'hf9a,
12'hf61,
12'hf36,
12'hf2c,
12'hf54,
12'hf97,
12'h001,
12'h084,
12'h0eb,
12'h100,
12'h0b5,
12'h04a,
12'hfee,
12'hfb8,
12'hfa9,
12'hfb6,
12'hfcd,
12'hfdf,
12'hffc,
12'h043,
12'h0df,
12'h1b8,
12'h26b,
12'h2a4,
12'h255,
12'h1d7,
12'h174,
12'h132,
12'h116,
12'h11b,
12'h140,
12'h17e,
12'h1bd,
12'h20e,
12'h286,
12'h2f8,
12'h324,
12'h2f4,
12'h28a,
12'h225,
12'h1e6,
12'h1d8,
12'h1f4,
12'h206,
12'h1ef,
12'h1ae,
12'h167,
12'h13b,
12'h125,
12'h125,
12'h133,
12'h142,
12'h142,
12'h127,
12'h100,
12'h0e9,
12'h0f3,
12'h0fe,
12'h0e4,
12'h0a1,
12'h053,
12'h00c,
12'hfd2,
12'hfad,
12'hf94,
12'hf7a,
12'hf4a,
12'heff,
12'hec9,
12'hedb,
12'hf28,
12'hf63,
12'hf70,
12'hf66,
12'hf52,
12'hf42,
12'hf3b,
12'hf4d,
12'hf5f,
12'hf42,
12'hef4,
12'he8e,
12'he66,
12'he87,
12'heb1,
12'hed7,
12'heea,
12'hee7,
12'hebf,
12'he6c,
12'he2c,
12'he3d,
12'he98,
12'hefe,
12'hf3a,
12'hf62,
12'hf91,
12'hf9a,
12'hf70,
12'hf4a,
12'hf4a,
12'hf60,
12'hf75,
12'hf90,
12'hfbb,
12'hfd9,
12'hfdb,
12'hfd5,
12'hfde,
12'hfe8,
12'hfda,
12'hfac,
12'hf7d,
12'hf84,
12'hfc0,
12'hffe,
12'h029,
12'h05d,
12'h0a3,
12'h0d7,
12'h0df,
12'h0c9,
12'h0c6,
12'h0ee,
12'h11b,
12'h130,
12'h11a,
12'h0ef,
12'h0bf,
12'h088,
12'h072,
12'h096,
12'h0ed,
12'h147,
12'h15c,
12'h12c,
12'h0e1,
12'h0bb,
12'h0b5,
12'h0ae,
12'h09b,
12'h082,
12'h067,
12'h048,
12'h03c,
12'h048,
12'h05f,
12'h080,
12'h08d,
12'h066,
12'h01c,
12'hfe2,
12'hfbd,
12'hfb1,
12'hfaa,
12'hf96,
12'hf89,
12'hf8b,
12'hf99,
12'hfa9,
12'hfb9,
12'hfbb,
12'hf96,
12'hf3c,
12'hecd,
12'he7d,
12'he5a,
12'he61,
12'he7c,
12'he9e,
12'hebb,
12'hec6,
12'hec7,
12'hebd,
12'hea7,
12'he82,
12'he5b,
12'he4d,
12'he5e,
12'he8f,
12'hedb,
12'hf2b,
12'hf5f,
12'hf60,
12'hf37,
12'hf13,
12'hefd,
12'hed5,
12'he9e,
12'he73,
12'he6c,
12'he83,
12'head,
12'hee9,
12'hf3f,
12'hfc5,
12'h057,
12'h0b2,
12'h0ae,
12'h060,
12'hff4,
12'hf87,
12'hf2c,
12'hee7,
12'hea7,
12'he74,
12'he64,
12'he8a,
12'hefe,
12'hfba,
12'h089,
12'h134,
12'h197,
12'h1a5,
12'h174,
12'h129,
12'h0d7,
12'h080,
12'h022,
12'hfd1,
12'hfa5,
12'hfc1,
12'h025,
12'h0b4,
12'h151,
12'h1e3,
12'h256,
12'h282,
12'h25d,
12'h20b,
12'h19b,
12'h10c,
12'h07e,
12'h049,
12'h0a6,
12'h17a,
12'h254,
12'h2ea,
12'h336,
12'h32e,
12'h2d9,
12'h257,
12'h1e8,
12'h1c6,
12'h1d0,
12'h1c0,
12'h17b,
12'h136,
12'h122,
12'h13d,
12'h16b,
12'h195,
12'h1a1,
12'h17e,
12'h128,
12'h0aa,
12'h03f,
12'h01c,
12'h039,
12'h055,
12'h04e,
12'h041,
12'h04d,
12'h073,
12'h086,
12'h066,
12'h012,
12'hf84,
12'hece,
12'he2c,
12'hde4,
12'he0d,
12'he72,
12'hed9,
12'hf1a,
12'hf35,
12'hf3c,
12'hf32,
12'hf20,
12'hf0f,
12'hefb,
12'heca,
12'he68,
12'hdf2,
12'hd98,
12'hd7b,
12'hda3,
12'he07,
12'he8b,
12'hf03,
12'hf35,
12'hf03,
12'he8f,
12'he21,
12'he17,
12'he80,
12'hf0b,
12'hf67,
12'hf82,
12'hf83,
12'hf7e,
12'hf6d,
12'hf5d,
12'hf60,
12'hf72,
12'hf7c,
12'hf77,
12'hf71,
12'hf82,
12'hfb0,
12'hfe6,
12'h010,
12'h02c,
12'h03d,
12'h041,
12'h039,
12'h02a,
12'h02a,
12'h050,
12'h094,
12'h0db,
12'h105,
12'h113,
12'h11c,
12'h137,
12'h16b,
12'h1ac,
12'h1f3,
12'h233,
12'h25a,
12'h25b,
12'h240,
12'h223,
12'h210,
12'h1ec,
12'h1ac,
12'h162,
12'h132,
12'h130,
12'h147,
12'h163,
12'h176,
12'h17f,
12'h173,
12'h13f,
12'h0f1,
12'h0b4,
12'h0b1,
12'h0d2,
12'h0ed,
12'h0ee,
12'h0db,
12'h0ca,
12'h0b0,
12'h090,
12'h078,
12'h060,
12'h03e,
12'h004,
12'hfcb,
12'hfaf,
12'hfb8,
12'hfcb,
12'hfc3,
12'hf9a,
12'hf56,
12'hf02,
12'heb0,
12'he77,
12'he57,
12'he3c,
12'he22,
12'he1c,
12'he3b,
12'he68,
12'he7b,
12'he6f,
12'he67,
12'he6e,
12'he5b,
12'he1e,
12'hde3,
12'hdd1,
12'hde4,
12'hdf9,
12'he05,
12'he27,
12'he65,
12'he8a,
12'he70,
12'he34,
12'he10,
12'he0b,
12'hdef,
12'hda6,
12'hd70,
12'hd90,
12'hdfd,
12'he6d,
12'heb1,
12'hed0,
12'hedb,
12'hec9,
12'he93,
12'he6c,
12'he83,
12'hec1,
12'hedf,
12'hec0,
12'heaf,
12'hef5,
12'hf81,
12'h00f,
12'h074,
12'h0ad,
12'h0b4,
12'h080,
12'h020,
12'hfbc,
12'hf7e,
12'hf73,
12'hf84,
12'hf97,
12'hfba,
12'h004,
12'h076,
12'h0fa,
12'h171,
12'h1c2,
12'h1ed,
12'h1eb,
12'h1c0,
12'h17f,
12'h138,
12'h0fb,
12'h0dc,
12'h0eb,
12'h134,
12'h1b3,
12'h262,
12'h317,
12'h396,
12'h3b1,
12'h362,
12'h2d4,
12'h24d,
12'h1fd,
12'h1e2,
12'h1e1,
12'h1e2,
12'h1e4,
12'h1e0,
12'h1d5,
12'h1cc,
12'h1ce,
12'h1d7,
12'h1d2,
12'h1ae,
12'h175,
12'h136,
12'h0fb,
12'h0c9,
12'h0ab,
12'h0a5,
12'h0b1,
12'h0be,
12'h0b7,
12'h096,
12'h068,
12'h03f,
12'h026,
12'h01b,
12'h007,
12'hfd1,
12'hf85,
12'hf49,
12'hf35,
12'hf3d,
12'hf42,
12'hf3d,
12'hf47,
12'hf6a,
12'hf9d,
12'hfc8,
12'hfdc,
12'hfcf,
12'hf93,
12'hf29,
12'hec1,
12'he97,
12'heb6,
12'hef0,
12'hf09,
12'hf00,
12'hef9,
12'hefd,
12'hef9,
12'hee3,
12'hed7,
12'hef2,
12'hf1f,
12'hf31,
12'hf25,
12'hf19,
12'hf15,
12'hf17,
12'hf1c,
12'hf36,
12'hf73,
12'hfb8,
12'hfd7,
12'hfd0,
12'hfc7,
12'hfd9,
12'h000,
12'h024,
12'h03a,
12'h038,
12'h014,
12'hfd8,
12'hfa6,
12'hf9f,
12'hfbc,
12'hfe0,
12'hfff,
12'h021,
12'h053,
12'h081,
12'h0af,
12'h0ea,
12'h132,
12'h16b,
12'h161,
12'h119,
12'h0cd,
12'h0a8,
12'h0a4,
12'h0a1,
12'h0a0,
12'h0ba,
12'h0dc,
12'h0e3,
12'h0d1,
12'h0c9,
12'h0d5,
12'h0cb,
12'h080,
12'h01a,
12'hff0,
12'h01f,
12'h074,
12'h0a7,
12'h0a8,
12'h099,
12'h08d,
12'h076,
12'h053,
12'h03d,
12'h041,
12'h045,
12'h032,
12'h016,
12'h018,
12'h03e,
12'h065,
12'h05b,
12'h016,
12'hfbb,
12'hf68,
12'hf1f,
12'hed3,
12'he92,
12'he84,
12'heb0,
12'hee9,
12'hef0,
12'hec0,
12'he84,
12'he62,
12'he62,
12'he78,
12'he9e,
12'hed2,
12'heff,
12'hefc,
12'hec0,
12'he75,
12'he59,
12'he74,
12'he94,
12'he9a,
12'he93,
12'he9d,
12'heb3,
12'heb5,
12'hea6,
12'hea6,
12'hec6,
12'hee5,
12'hed7,
12'he9b,
12'he64,
12'he5c,
12'he8e,
12'hedd,
12'hf2b,
12'hf58,
12'hf4c,
12'hef5,
12'he6d,
12'he00,
12'hde8,
12'he2c,
12'he9a,
12'hf01,
12'hf61,
12'hfcf,
12'h04e,
12'h0d2,
12'h13b,
12'h171,
12'h15c,
12'h0f0,
12'h045,
12'hf96,
12'hf26,
12'hf27,
12'hf94,
12'h02c,
12'h0b4,
12'h110,
12'h153,
12'h1a2,
12'h20f,
12'h27b,
12'h2ae,
12'h280,
12'h1fa,
12'h154,
12'h0c9,
12'h09b,
12'h0ef,
12'h1b2,
12'h288,
12'h30e,
12'h32b,
12'h313,
12'h2f8,
12'h2d5,
12'h2a1,
12'h269,
12'h247,
12'h229,
12'h1ea,
12'h18d,
12'h156,
12'h175,
12'h1c5,
12'h203,
12'h207,
12'h1d7,
12'h178,
12'h0ec,
12'h053,
12'hff7,
12'h006,
12'h057,
12'h08c,
12'h084,
12'h06b,
12'h06f,
12'h08b,
12'h09b,
12'h084,
12'h036,
12'hfb6,
12'hf13,
12'he89,
12'he5c,
12'he99,
12'hf0c,
12'hf74,
12'hfad,
12'hfb5,
12'hf99,
12'hf6b,
12'hf3b,
12'hf09,
12'heb7,
12'he37,
12'hda8,
12'hd43,
12'hd35,
12'hd7d,
12'he07,
12'heba,
12'hf61,
12'hfbf,
12'hfb9,
12'hf78,
12'hf40,
12'hf2e,
12'hf2e,
12'hf22,
12'hefe,
12'heca,
12'he8c,
12'he56,
12'he41,
12'he57,
12'he94,
12'hee4,
12'hf3f,
12'hfa6,
12'h015,
12'h079,
12'h0bc,
12'h0cf,
12'h0ac,
12'h056,
12'hfe5,
12'hf7c,
12'hf31,
12'hf0a,
12'hf0f,
12'hf55,
12'hfdc,
12'h07d,
12'h106,
12'h163,
12'h1a2,
12'h1c6,
12'h1be,
12'h18d,
12'h15c,
12'h15c,
12'h18c,
12'h1c0,
12'h1d3,
12'h1ca,
12'h1bb,
12'h1a9,
12'h18f,
12'h17b,
12'h183,
12'h196,
12'h18c,
12'h153,
12'h10c,
12'h0ef,
12'h10c,
12'h136,
12'h12f,
12'h0f0,
12'h0a4,
12'h076,
12'h073,
12'h08a,
12'h0ae,
12'h0d7,
12'h0f1,
12'h0dd,
12'h094,
12'h03c,
12'h003,
12'hfe7,
12'hfcc,
12'hfa9,
12'hf90,
12'hf91,
12'hf8f,
12'hf60,
12'hf04,
12'hea5,
12'he65,
12'he41,
12'he2a,
12'he24,
12'he37,
12'he58,
12'he6c,
12'he6d,
12'he6d,
12'he79,
12'he8c,
12'he9a,
12'he91,
12'he66,
12'he1b,
12'hdce,
12'hda6,
12'hdb4,
12'hdee,
12'he45,
12'hea3,
12'hee9,
12'hef1,
12'heb9,
12'he7e,
12'he7b,
12'heae,
12'hee0,
12'hef3,
12'hef4,
12'hef0,
12'hed6,
12'he9b,
12'he6c,
12'he80,
12'hed5,
12'hf24,
12'hf35,
12'hf1f,
12'hf16,
12'hf21,
12'hf36,
12'hf64,
12'hfc8,
12'h055,
12'h0d1,
12'h110,
12'h116,
12'h0fa,
12'h0c2,
12'h066,
12'hfef,
12'hf7d,
12'hf38,
12'hf34,
12'hf6d,
12'hfcf,
12'h042,
12'h0bc,
12'h13c,
12'h1b5,
12'h20e,
12'h22a,
12'h207,
12'h1bd,
12'h15c,
12'h0ec,
12'h08a,
12'h06f,
12'h0c1,
12'h156,
12'h1ea,
12'h25f,
12'h2bc,
12'h2f7,
12'h2e4,
12'h281,
12'h209,
12'h1c6,
12'h1bd,
12'h1b9,
12'h19f,
12'h17f,
12'h167,
12'h14f,
12'h135,
12'h12a,
12'h13c,
12'h150,
12'h141,
12'h109,
12'h0ca,
12'h0a7,
12'h0ab,
12'h0c6,
12'h0e0,
12'h0e9,
12'h0d0,
12'h097,
12'h05b,
12'h03b,
12'h035,
12'h034,
12'h025,
12'hff2,
12'hf8c,
12'hf11,
12'hec1,
12'hed4,
12'hf3f,
12'hfb7,
12'hff8,
12'hff1,
12'hfaf,
12'hf4b,
12'hef2,
12'hed5,
12'hf00,
12'hf43,
12'hf51,
12'hf0e,
12'hea0,
12'he4c,
12'he47,
12'he95,
12'hf12,
12'hf89,
12'hfb8,
12'hf85,
12'hf1c,
12'hec4,
12'heb1,
12'hee4,
12'hf39,
12'hf74,
12'hf61,
12'hf05,
12'he9d,
12'he70,
12'he9b,
12'heff,
12'hf6c,
12'hfc6,
12'h003,
12'h01f,
12'h029,
12'h046,
12'h087,
12'h0bb,
12'h09b,
12'h020,
12'hf88,
12'hf25,
12'hf1b,
12'hf59,
12'hfbe,
12'h02f,
12'h084,
12'h096,
12'h077,
12'h066,
12'h08f,
12'h0e8,
12'h13f,
12'h168,
12'h151,
12'h108,
12'h0b1,
12'h078,
12'h075,
12'h09d,
12'h0c8,
12'h0da,
12'h0ca,
12'h09d,
12'h065,
12'h047,
12'h061,
12'h0a0,
12'h0cd,
12'h0c3,
12'h095,
12'h070,
12'h064,
12'h062,
12'h067,
12'h078,
12'h083,
12'h069,
12'h01e,
12'hfd3,
12'hfb7,
12'hfc4,
12'hfce,
12'hfc2,
12'hfad,
12'hfa1,
12'hf9e,
12'hfa6,
12'hfbf,
12'hfe2,
12'hff0,
12'hfcc,
12'hf7f,
12'hf29,
12'heee,
12'hed9,
12'hee1,
12'hef1,
12'hef7,
12'heee,
12'hedf,
12'hedd,
12'hef0,
12'hf02,
12'hf02,
12'hef8,
12'hef4,
12'hef8,
12'hf06,
12'hf36,
12'hf8a,
12'hfd8,
12'hfea,
12'hfaa,
12'hf3e,
12'hed6,
12'he85,
12'he4f,
12'he3d,
12'he56,
12'he84,
12'he98,
12'he86,
12'he7e,
12'heb0,
12'hf18,
12'hf8f,
12'hfe5,
12'h000,
12'hfd7,
12'hf69,
12'hed8,
12'he61,
12'he39,
12'he65,
12'heba,
12'hf14,
12'hf65,
12'hfb2,
12'h016,
12'h09f,
12'h136,
12'h1a2,
12'h1aa,
12'h14c,
12'h0a4,
12'hfdb,
12'hf2d,
12'hecd,
12'hede,
12'hf46,
12'hfd3,
12'h064,
12'h107,
12'h1d0,
12'h2a4,
12'h348,
12'h385,
12'h343,
12'h28e,
12'h18d,
12'h092,
12'h00c,
12'h03b,
12'h0f9,
12'h1cf,
12'h25c,
12'h290,
12'h287,
12'h270,
12'h276,
12'h29f,
12'h2cf,
12'h2cd,
12'h26f,
12'h1c2,
12'h10a,
12'h09c,
12'h099,
12'h0ee,
12'h15f,
12'h1a3,
12'h19c,
12'h15d,
12'h11e,
12'h0fe,
12'h0f4,
12'h0f9,
12'h0fa,
12'h0ec,
12'h0d0,
12'h0b3,
12'h0b4,
12'h0da,
12'h0f8,
12'h0c0,
12'h020,
12'hf51,
12'he9e,
12'he3d,
12'he47,
12'hea9,
12'hf24,
12'hf71,
12'hf74,
12'hf55,
12'hf5e,
12'hfb0,
12'h01c,
12'h056,
12'h019,
12'hf68,
12'he69,
12'hd7b,
12'hd06,
12'hd33,
12'hddc,
12'hea3,
12'hf3a,
12'hf7e,
12'hf71,
12'hf29,
12'hedb,
12'hebb,
12'hed6,
12'hef7,
12'hef2,
12'hed0,
12'heab,
12'he92,
12'he8f,
12'hea4,
12'hed4,
12'hf0a,
12'hf2f,
12'hf40,
12'hf54,
12'hf7e,
12'hfa5,
12'hfb2,
12'hfa4,
12'hf99,
12'hf95,
12'hf90,
12'hf91,
12'hfa7,
12'hfd3,
12'hff8,
12'h000,
12'hffc,
12'h00c,
12'h03d,
12'h084,
12'h0d0,
12'h119,
12'h15e,
12'h190,
12'h19f,
12'h198,
12'h193,
12'h19f,
12'h1b5,
12'h1b5,
12'h18c,
12'h141,
12'h0fe,
12'h0d7,
12'h0d7,
12'h102,
12'h132,
12'h155,
12'h160,
12'h150,
12'h12c,
12'h108,
12'h100,
12'h109,
12'h101,
12'h0d2,
12'h090,
12'h05e,
12'h051,
12'h061,
12'h075,
12'h068,
12'h041,
12'h00c,
12'hfdc,
12'hfc9,
12'hfd7,
12'hff5,
12'h007,
12'hff9,
12'hfa8,
12'hf23,
12'he8f,
12'he21,
12'hdfc,
12'he17,
12'he4d,
12'he77,
12'he93,
12'hea9,
12'heca,
12'hef1,
12'hf0f,
12'hf0c,
12'hed4,
12'he7b,
12'he20,
12'hde3,
12'hdce,
12'hde8,
12'he2a,
12'he85,
12'hee4,
12'hf1a,
12'hf2b,
12'hf2a,
12'hf1e,
12'hef4,
12'he99,
12'he3d,
12'he0b,
12'he0e,
12'he34,
12'he60,
12'he83,
12'he97,
12'hea9,
12'hec4,
12'heea,
12'hf13,
12'hf1f,
12'hefb,
12'hec3,
12'hea4,
12'hec9,
12'hf45,
12'hff8,
12'h0aa,
12'h119,
12'h119,
12'h0c4,
12'h05c,
12'h00e,
12'hfd0,
12'hf86,
12'hf3f,
12'hf05,
12'heea,
12'hf0f,
12'hf9c,
12'h0a4,
12'h1cc,
12'h293,
12'h2a7,
12'h231,
12'h1a6,
12'h146,
12'h11a,
12'h100,
12'h0e8,
12'h0db,
12'h0ee,
12'h136,
12'h1ca,
12'h29e,
12'h363,
12'h3bd,
12'h384,
12'h2eb,
12'h244,
12'h1e7,
12'h1ff,
12'h266,
12'h2af,
12'h279,
12'h1e2,
12'h15f,
12'h146,
12'h192,
12'h209,
12'h258,
12'h256,
12'h1f4,
12'h147,
12'h0ad,
12'h094,
12'h101,
12'h18e,
12'h1c3,
12'h184,
12'h107,
12'h08f,
12'h046,
12'h037,
12'h056,
12'h06a,
12'h037,
12'hfc3,
12'hf57,
12'hf53,
12'hfa9,
12'hff4,
12'h004,
12'hfd8,
12'hf6f,
12'hee1,
12'he61,
12'he41,
12'he89,
12'hef2,
12'hf28,
12'hf0c,
12'hed0,
12'head,
12'heac,
12'hebc,
12'hed1,
12'hed5,
12'heb8,
12'he8a,
12'he62,
12'he54,
12'he6a,
12'hea6,
12'hef1,
12'hf28,
12'hf3c,
12'hf23,
12'hef3,
12'hed0,
12'hece,
12'hedf,
12'hef9,
12'hf32,
12'hf85,
12'hfd5,
12'hffc,
12'hffb,
12'hfe4,
12'hfce,
12'hfb7,
12'hf87,
12'hf57,
12'hf3f,
12'hf4e,
12'hf6f,
12'hf96,
12'hfda,
12'h038,
12'h0aa,
12'h100,
12'h124,
12'h123,
12'h122,
12'h136,
12'h145,
12'h140,
12'h112,
12'h0c5,
12'h082,
12'h072,
12'h09a,
12'h0d5,
12'h10f,
12'h130,
12'h118,
12'h0cd,
12'h081,
12'h06c,
12'h08c,
12'h0b7,
12'h0b5,
12'h07b,
12'h044,
12'h044,
12'h06f,
12'h0a3,
12'h0c6,
12'h0b9,
12'h062,
12'hfe2,
12'hf7f,
12'hf60,
12'hf8b,
12'hfe9,
12'h042,
12'h05c,
12'h02c,
12'hfe6,
12'hfc9,
12'hfe5,
12'hffb,
12'hfd5,
12'hf64,
12'hebc,
12'he10,
12'hd96,
12'hd8e,
12'he03,
12'heac,
12'hf42,
12'hf92,
12'hf81,
12'hf34,
12'hee3,
12'hec0,
12'hec5,
12'hed4,
12'hee9,
12'hedc,
12'heaf,
12'he83,
12'he8a,
12'hed9,
12'hf2e,
12'hf5a,
12'hf58,
12'hf4f,
12'hf54,
12'hf53,
12'hf51,
12'hf49,
12'hf33,
12'hf09,
12'hec8,
12'he95,
12'he8d,
12'head,
12'heea,
12'hf22,
12'hf44,
12'hf4d,
12'hf30,
12'hef4,
12'heaa,
12'he60,
12'he25,
12'he17,
12'he44,
12'he9d,
12'hf0c,
12'hf7f,
12'h000,
12'h08c,
12'h104,
12'h14e,
12'h14c,
12'h102,
12'h07e,
12'hfe1,
12'hf5c,
12'hf14,
12'hf29,
12'hf97,
12'h029,
12'h0c4,
12'h150,
12'h1c2,
12'h226,
12'h279,
12'h2bc,
12'h2cb,
12'h28d,
12'h1e5,
12'h0e0,
12'h01d,
12'h014,
12'h0ca,
12'h1e8,
12'h2f9,
12'h3b6,
12'h3ff,
12'h3eb,
12'h3a9,
12'h357,
12'h315,
12'h2cd,
12'h24d,
12'h1a0,
12'h0fc,
12'h098,
12'h096,
12'h0fd,
12'h1a3,
12'h23d,
12'h292,
12'h292,
12'h23f,
12'h1b6,
12'h138,
12'h0e2,
12'h088,
12'h012,
12'hfa0,
12'hf76,
12'hfac,
12'h013,
12'h09b,
12'h106,
12'h12b,
12'h0fa,
12'h068,
12'hfb9,
12'hf2e,
12'hede,
12'hebf,
12'heac,
12'he99,
12'he8b,
12'he8e,
12'hec7,
12'hf2d,
12'hf80,
12'hf81,
12'hf22,
12'he93,
12'he13,
12'hdbe,
12'hda5,
12'hdc4,
12'he02,
12'he44,
12'he6d,
12'he80,
12'he90,
12'he9c,
12'he9e,
12'he96,
12'he9f,
12'hec5,
12'heed,
12'hefa,
12'hedd,
12'heaa,
12'he6b,
12'he3c,
12'he40,
12'he99,
12'hf3f,
12'hfe4,
12'h044,
12'h052,
12'h02a,
12'hff8,
12'hfcb,
12'hf9c,
12'hf7b,
12'hf70,
12'hf84,
12'hf9a,
12'hfac,
12'hff1,
12'h06b,
12'h0ed,
12'h140,
12'h15b,
12'h159,
12'h152,
12'h167,
12'h184,
12'h1a1,
12'h1cd,
12'h1de,
12'h1ce,
12'h1a0,
12'h162,
12'h138,
12'h130,
12'h148,
12'h178,
12'h1ad,
12'h1c3,
12'h19b,
12'h145,
12'h0ee,
12'h0ba,
12'h0b5,
12'h0ca,
12'h0e9,
12'h103,
12'h11c,
12'h136,
12'h152,
12'h163,
12'h162,
12'h14f,
12'h118,
12'h0b8,
12'h031,
12'hfb2,
12'hf6a,
12'hf5d,
12'hf92,
12'hfe8,
12'h01f,
12'h02b,
12'h006,
12'hfb2,
12'hf3b,
12'heae,
12'he22,
12'hdcd,
12'hdb0,
12'hda4,
12'hd97,
12'hda0,
12'hde6,
12'he50,
12'hea5,
12'heb3,
12'he93,
12'he59,
12'hdee,
12'hd7a,
12'hd51,
12'hd76,
12'hdb3,
12'hde3,
12'he09,
12'he4d,
12'he97,
12'hea4,
12'he81,
12'he66,
12'he6c,
12'he73,
12'he5c,
12'he43,
12'he4c,
12'he77,
12'he8b,
12'he75,
12'he5f,
12'he7f,
12'hedd,
12'hf2d,
12'hf42,
12'hf40,
12'hf33,
12'hf18,
12'hf05,
12'hf1e,
12'hf75,
12'hfbb,
12'hfbb,
12'hfb6,
12'h00d,
12'h0bb,
12'h151,
12'h16e,
12'h103,
12'h045,
12'hf91,
12'hf2f,
12'hf47,
12'hfd4,
12'h07b,
12'h100,
12'h165,
12'h1cc,
12'h22d,
12'h276,
12'h290,
12'h273,
12'h22e,
12'h1bb,
12'h142,
12'h100,
12'h129,
12'h1d0,
12'h299,
12'h329,
12'h380,
12'h3ab,
12'h3c0,
12'h3aa,
12'h36d,
12'h329,
12'h2ca,
12'h262,
12'h212,
12'h1f1,
12'h200,
12'h219,
12'h227,
12'h21c,
12'h1fd,
12'h1d2,
12'h19d,
12'h190,
12'h1a9,
12'h1be,
12'h1ad,
12'h165,
12'h0fa,
12'h095,
12'h058,
12'h040,
12'h04d,
12'h064,
12'h053,
12'h013,
12'hfbe,
12'hf91,
12'hfa5,
12'hfa8,
12'hf65,
12'hef9,
12'hea4,
12'he9a,
12'hec5,
12'hefa,
12'hf23,
12'hf23,
12'heef,
12'hea8,
12'he86,
12'hea0,
12'hecf,
12'hed6,
12'hea0,
12'he56,
12'he16,
12'hdfd,
12'he12,
12'he4b,
12'he8a,
12'hea9,
12'he93,
12'he68,
12'he71,
12'hebb,
12'hf08,
12'hf24,
12'hf09,
12'hed1,
12'he8f,
12'he4d,
12'he36,
12'he7a,
12'hef0,
12'hf53,
12'hf98,
12'hfaf,
12'hfc4,
12'hfeb,
12'hffa,
12'hffc,
12'hff7,
12'hfcd,
12'hf68,
12'hf03,
12'hef2,
12'hf51,
12'hfea,
12'h06a,
12'h0c9,
12'h103,
12'h10e,
12'h0f0,
12'h0bd,
12'h0b3,
12'h0ee,
12'h121,
12'h118,
12'h0f0,
12'h0e1,
12'h105,
12'h130,
12'h146,
12'h14a,
12'h130,
12'h108,
12'h0dd,
12'h0c1,
12'h0b9,
12'h0be,
12'h0d2,
12'h0d6,
12'h0c8,
12'h0b2,
12'h0a7,
12'h0b5,
12'h0b3,
12'h097,
12'h086,
12'h0a1,
12'h0c9,
12'h0c6,
12'h093,
12'h055,
12'h01d,
12'hfe7,
12'hfb7,
12'hfa2,
12'hfc1,
12'hfe3,
12'hfda,
12'hfc0,
12'hfa2,
12'hf7f,
12'hf48,
12'hf17,
12'hf08,
12'hef8,
12'heda,
12'heb4,
12'he97,
12'hea1,
12'hec0,
12'hed5,
12'hee3,
12'hee7,
12'hec8,
12'he9b,
12'he71,
12'he67,
12'he93,
12'hec5,
12'hefa,
12'hf1b,
12'hf15,
12'hefa,
12'hecc,
12'hebb,
12'hec4,
12'heaf,
12'he6e,
12'he2c,
12'he1a,
12'he30,
12'he42,
12'he41,
12'he5c,
12'heb5,
12'hf25,
12'hf61,
12'hf70,
12'hf6c,
12'hf57,
12'hf3e,
12'hf21,
12'hefb,
12'hed8,
12'hebf,
12'hea5,
12'he9d,
12'hec1,
12'hf19,
12'hf9e,
12'h043,
12'h0f4,
12'h16b,
12'h18a,
12'h164,
12'h104,
12'h07c,
12'hfdb,
12'hf57,
12'hf29,
12'hf4a,
12'hfad,
12'h04c,
12'h11a,
12'h1fd,
12'h2b8,
12'h30e,
12'h31a,
12'h2f5,
12'h292,
12'h1e2,
12'h111,
12'h08d,
12'h0a1,
12'h154,
12'h241,
12'h304,
12'h378,
12'h392,
12'h378,
12'h348,
12'h319,
12'h2ef,
12'h2b7,
12'h270,
12'h227,
12'h1db,
12'h180,
12'h137,
12'h140,
12'h198,
12'h1f0,
12'h209,
12'h1e5,
12'h1ae,
12'h180,
12'h15d,
12'h149,
12'h131,
12'h0fd,
12'h0b6,
12'h06f,
12'h031,
12'h017,
12'h020,
12'h036,
12'h037,
12'hfed,
12'hf52,
12'heb9,
12'he70,
12'he81,
12'hec0,
12'hedf,
12'hebb,
12'he73,
12'he49,
12'he77,
12'heea,
12'hf54,
12'hf6f,
12'hf10,
12'he4a,
12'hd85,
12'hd1a,
12'hd2f,
12'hdb2,
12'he5a,
12'hee6,
12'hf26,
12'hf10,
12'hec6,
12'he70,
12'he43,
12'he56,
12'he80,
12'he87,
12'he74,
12'he5c,
12'he47,
12'he63,
12'heb6,
12'hf12,
12'hf57,
12'hf83,
12'hf96,
12'hf9c,
12'hfa9,
12'hfce,
12'h010,
12'h04a,
12'h064,
12'h058,
12'h014,
12'hfbd,
12'hf74,
12'hf6a,
12'hfaa,
12'h002,
12'h05a,
12'h0b0,
12'h102,
12'h14c,
12'h17d,
12'h191,
12'h1a9,
12'h1cc,
12'h1da,
12'h1c9,
12'h1a5,
12'h18d,
12'h187,
12'h17d,
12'h17c,
12'h18b,
12'h1a6,
12'h1b1,
12'h188,
12'h14c,
12'h10c,
12'h0e9,
12'h109,
12'h154,
12'h18e,
12'h187,
12'h145,
12'h0f2,
12'h0d3,
12'h0f1,
12'h11e,
12'h135,
12'h11f,
12'h0e3,
12'h092,
12'h03c,
12'h00c,
12'h021,
12'h043,
12'h03f,
12'h018,
12'hfd0,
12'hf75,
12'hf37,
12'hf19,
12'heff,
12'hec1,
12'he59,
12'he07,
12'hde5,
12'hde7,
12'he06,
12'he29,
12'he3a,
12'he4a,
12'he61,
12'he77,
12'he76,
12'he54,
12'he24,
12'hdf0,
12'hdc9,
12'hda4,
12'hd79,
12'hd7c,
12'hdda,
12'he69,
12'hee7,
12'hf27,
12'hf17,
12'heef,
12'heb9,
12'he57,
12'hdea,
12'hdba,
12'hde3,
12'he2b,
12'he6b,
12'he8f,
12'he98,
12'heb6,
12'hee2,
12'hf0b,
12'hf1e,
12'hf10,
12'hefa,
12'hed6,
12'heb9,
12'hee6,
12'hf81,
12'h046,
12'h0ea,
12'h143,
12'h14c,
12'h114,
12'h096,
12'h010,
12'hfb6,
12'hf88,
12'hf74,
12'hf79,
12'hfa8,
12'hfee,
12'h050,
12'h0ee,
12'h1b2,
12'h249,
12'h262,
12'h1fa,
12'h175,
12'h143,
12'h15b,
12'h163,
12'h146,
12'h138,
12'h16c,
12'h1d9,
12'h25e,
12'h2f1,
12'h392,
12'h3f9,
12'h3d7,
12'h33a,
12'h298,
12'h244,
12'h227,
12'h234,
12'h24e,
12'h23f,
12'h1fd,
12'h1c0,
12'h1cd,
12'h21a,
12'h25d,
12'h255,
12'h201,
12'h180,
12'h0f3,
12'h07e,
12'h053,
12'h097,
12'h0f0,
12'h10c,
12'h102,
12'h0df,
12'h0b1,
12'h07f,
12'h055,
12'h046,
12'h02d,
12'hfdf,
12'hf52,
12'hec8,
12'he8c,
12'he9e,
12'hec7,
12'hedc,
12'heec,
12'hefd,
12'hef9,
12'hecf,
12'he9f,
12'he99,
12'heaf,
12'heb1,
12'he99,
12'he7f,
12'he71,
12'he7c,
12'he99,
12'heb1,
12'heaa,
12'he9d,
12'he95,
12'he8c,
12'he88,
12'he83,
12'he94,
12'hebb,
12'heed,
12'hf21,
12'hf39,
12'hf25,
12'hefe,
12'hee1,
12'hee3,
12'hf10,
12'hf72,
12'hfef,
12'h040,
12'h03d,
12'h004,
12'hfc6,
12'hfa8,
12'hfae,
12'hfbf,
12'hfce,
12'hfc5,
12'hfaa,
12'hf9d,
12'hfa2,
12'hfd2,
12'h052,
12'h0f1,
12'h150,
12'h14a,
12'h110,
12'h0eb,
12'h0fa,
12'h136,
12'h16f,
12'h185,
12'h165,
12'h11b,
12'h0da,
12'h0bc,
12'h0cf,
12'h10c,
12'h155,
12'h17a,
12'h14e,
12'h0e0,
12'h08e,
12'h081,
12'h09d,
12'h0c0,
12'h0c4,
12'h0bc,
12'h0b7,
12'h0aa,
12'h090,
12'h075,
12'h066,
12'h061,
12'h03d,
12'hfed,
12'hfa1,
12'hf8d,
12'hfba,
12'hff6,
12'h017,
12'h01d,
12'h00b,
12'hfe3,
12'hfb9,
12'hfa5,
12'hf8c,
12'hf44,
12'hec5,
12'he31,
12'hdd5,
12'hdc3,
12'hdec,
12'he50,
12'heb4,
12'hef5,
12'hef9,
12'hed6,
12'hec0,
12'heab,
12'he93,
12'he76,
12'he6e,
12'he9c,
12'hec2,
12'heac,
12'he86,
12'he9f,
12'hefb,
12'hf2f,
12'hf1e,
12'hf02,
12'hf03,
12'hf26,
12'hf34,
12'hf22,
12'hf31,
12'hf4c,
12'hf2e,
12'hee4,
12'hea4,
12'heb2,
12'heff,
12'hf45,
12'hf83,
12'hfd5,
12'h01a,
12'h017,
12'hfb0,
12'hf37,
12'hee7,
12'hea5,
12'he7e,
12'he77,
12'hea7,
12'hf0f,
12'hf95,
12'h041,
12'h100,
12'h1b9,
12'h21f,
12'h210,
12'h1ab,
12'h0fd,
12'h028,
12'hf71,
12'hf18,
12'hf2a,
12'hf94,
12'h01b,
12'h088,
12'h0df,
12'h142,
12'h1c5,
12'h25a,
12'h2d8,
12'h315,
12'h2d0,
12'h204,
12'h109,
12'h058,
12'h060,
12'h107,
12'h1d3,
12'h26f,
12'h2d1,
12'h312,
12'h339,
12'h34c,
12'h346,
12'h30c,
12'h299,
12'h1ef,
12'h12a,
12'h090,
12'h05d,
12'h094,
12'h103,
12'h17b,
12'h1d2,
12'h1fb,
12'h1fa,
12'h1ce,
12'h180,
12'h135,
12'h0f4,
12'h0ab,
12'h045,
12'hfce,
12'hf96,
12'hfbe,
12'h011,
12'h049,
12'h043,
12'hff4,
12'hf71,
12'hef5,
12'heac,
12'heb7,
12'hefd,
12'hf34,
12'hf33,
12'hf05,
12'hec4,
12'hea9,
12'hed2,
12'hf13,
12'hf36,
12'hf0d,
12'he9d,
12'he12,
12'hd95,
12'hd61,
12'hd82,
12'hde3,
12'he64,
12'heb9,
12'hed0,
12'hebe,
12'heb5,
12'hee0,
12'hf29,
12'hf6d,
12'hf79,
12'hf4c,
12'hef8,
12'he96,
12'he45,
12'he20,
12'he47,
12'he9d,
12'hf07,
12'hf6f,
12'hfc5,
12'h010,
12'h049,
12'h066,
12'h07a,
12'h08d,
12'h070,
12'h018,
12'hfbe,
12'hf8e,
12'hfa3,
12'hff3,
12'h05b,
12'h0b3,
12'h0ee,
12'h108,
12'h105,
12'h10c,
12'h127,
12'h156,
12'h190,
12'h1c5,
12'h1f0,
12'h1f9,
12'h1de,
12'h1bc,
12'h191,
12'h16e,
12'h167,
12'h165,
12'h174,
12'h18d,
12'h194,
12'h17e,
12'h147,
12'h119,
12'h111,
12'h114,
12'h0f3,
12'h0b8,
12'h09e,
12'h0b9,
12'h0e9,
12'h10a,
12'h109,
12'h106,
12'h0ff,
12'h0c4,
12'h062,
12'h00a,
12'hfd7,
12'hfba,
12'hf9f,
12'hfa4,
12'hfce,
12'h002,
12'h01b,
12'hffd,
12'hfb4,
12'hf3d,
12'heaa,
12'he22,
12'hdc3,
12'hd96,
12'hd87,
12'hda1,
12'hde5,
12'he36,
12'he77,
12'hea3,
12'hec5,
12'hec5,
12'he92,
12'he3a,
12'hde9,
12'hdc1,
12'hdb0,
12'hd9c,
12'hda0,
12'hde5,
12'he4f,
12'hea4,
12'heca,
12'hec4,
12'heca,
12'hee3,
12'hed0,
12'he83,
12'he21,
12'hdea,
12'hde9,
12'he20,
12'he7e,
12'hedc,
12'hf2f,
12'hf4e,
12'hf2c,
12'hf04,
12'hef9,
12'hf05,
12'hf19,
12'hf1d,
12'hf18,
12'hf30,
12'hf6f,
12'hfdc,
12'h080,
12'h12f,
12'h1a0,
12'h189,
12'h0f8,
12'h04a,
12'hfb9,
12'hf66,
12'hf51,
12'hf72,
12'hfa1,
12'hfcf,
12'h037,
12'h0e8,
12'h1b3,
12'h23f,
12'h258,
12'h22d,
12'h1ea,
12'h194,
12'h147,
12'h130,
12'h160,
12'h1c8,
12'h223,
12'h24f,
12'h26a,
12'h292,
12'h2d4,
12'h2eb,
12'h2c1,
12'h286,
12'h25b,
12'h24b,
12'h268,
12'h2aa,
12'h2c4,
12'h28b,
12'h217,
12'h1b2,
12'h180,
12'h15f,
12'h140,
12'h11f,
12'h108,
12'h0fa,
12'h0fc,
12'h102,
12'h116,
12'h144,
12'h157,
12'h146,
12'h0ff,
12'h097,
12'h024,
12'hfbc,
12'hf85,
12'hf6c,
12'hf56,
12'hf28,
12'heec,
12'hecb,
12'heeb,
12'hf44,
12'hf91,
12'hfc0,
12'hfd5,
12'hfab,
12'hf56,
12'hf05,
12'hecf,
12'hebc,
12'hea3,
12'he68,
12'he40,
12'he47,
12'he81,
12'hed3,
12'hf14,
12'hf29,
12'hf05,
12'heb6,
12'he5f,
12'he4f,
12'he95,
12'hef3,
12'hf40,
12'hf7c,
12'hf99,
12'hf96,
12'hf6b,
12'hf24,
12'hefc,
12'hf05,
12'hf1e,
12'hf23,
12'hf3c,
12'hf8c,
12'hff7,
12'h04a,
12'h061,
12'h03e,
12'hffe,
12'hfb0,
12'hf78,
12'hf6c,
12'hf86,
12'hfbe,
12'hfe0,
12'hfd4,
12'hfe4,
12'h02b,
12'h0a1,
12'h11e,
12'h162,
12'h16e,
12'h14d,
12'h116,
12'h0ee,
12'h0ea,
12'h0f3,
12'h0f3,
12'h0e9,
12'h0e0,
12'h0e4,
12'h0eb,
12'h0ff,
12'h114,
12'h10e,
12'h0e0,
12'h08f,
12'h04b,
12'h034,
12'h03b,
12'h04a,
12'h060,
12'h07b,
12'h08b,
12'h08b,
12'h08d,
12'h097,
12'h093,
12'h068,
12'h013,
12'hfb9,
12'hf80,
12'hf78,
12'hf9a,
12'hfd4,
12'h015,
12'h033,
12'h015,
12'hfc2,
12'hf5a,
12'hf01,
12'hec6,
12'he94,
12'he67,
12'he49,
12'he39,
12'he4c,
12'he86,
12'hed7,
12'hf07,
12'hef5,
12'hebe,
12'he8a,
12'he7a,
12'he7f,
12'he8e,
12'hebe,
12'hf06,
12'hf31,
12'hf30,
12'hf2d,
12'hf4c,
12'hf6e,
12'hf5d,
12'hf27,
12'hf05,
12'hf0f,
12'hf20,
12'hf1a,
12'hf2d,
12'hf5b,
12'hf83,
12'hf7e,
12'hf40,
12'hf07,
12'hf10,
12'hf64,
12'hfc2,
12'hfe7,
12'hfbd,
12'hf57,
12'hee4,
12'he97,
12'he6d,
12'he5c,
12'he5c,
12'he6e,
12'heab,
12'hf20,
12'hfd9,
12'h0a9,
12'h177,
12'h20d,
12'h223,
12'h1ab,
12'h0d9,
12'h014,
12'hf73,
12'hef7,
12'hec3,
12'hedb,
12'hf47,
12'hfdc,
12'h073,
12'h129,
12'h1ed,
12'h284,
12'h2dc,
12'h2e2,
12'h28f,
12'h1f7,
12'h11f,
12'h059,
12'hff5,
12'h008,
12'h0ac,
12'h19d,
12'h27b,
12'h313,
12'h358,
12'h365,
12'h35b,
12'h33f,
12'h300,
12'h296,
12'h214,
12'h1a3,
12'h14b,
12'h0ec,
12'h099,
12'h08e,
12'h0ed,
12'h189,
12'h215,
12'h26a,
12'h262,
12'h1eb,
12'h134,
12'h08a,
12'h02d,
12'h00b,
12'h012,
12'h03a,
12'h04f,
12'h046,
12'h038,
12'h03b,
12'h051,
12'h051,
12'h01c,
12'hfb1,
12'hf37,
12'heef,
12'hef4,
12'hf38,
12'hf6a,
12'hf42,
12'hef0,
12'heba,
12'hea8,
12'he9e,
12'he9b,
12'hea5,
12'hea6,
12'he83,
12'he43,
12'he11,
12'he13,
12'he50,
12'heb1,
12'hf0f,
12'hf4a,
12'hf4c,
12'hf09,
12'heb6,
12'he9b,
12'hecb,
12'hf21,
12'hf5d,
12'hf4e,
12'hefe,
12'hea1,
12'he6e,
12'he6b,
12'he95,
12'hee4,
12'hf45,
12'hfaa,
12'hff9,
12'h01e,
12'h029,
12'h023,
12'h019,
12'h009,
12'hfe1,
12'hfa9,
12'hf8f,
12'hf9f,
12'hfb5,
12'hfd3,
12'h003,
12'h03f,
12'h07e,
12'h0b1,
12'h0d6,
12'h0fa,
12'h11f,
12'h150,
12'h185,
12'h1b8,
12'h1d1,
12'h1af,
12'h166,
12'h113,
12'h0d5,
12'h0c1,
12'h0db,
12'h103,
12'h119,
12'h113,
12'h0db,
12'h07f,
12'h034,
12'h021,
12'h058,
12'h0b4,
12'h0e9,
12'h0ea,
12'h0bf,
12'h08a,
12'h079,
12'h098,
12'h0dc,
12'h101,
12'h0dc,
12'h05f,
12'hfbb,
12'hf53,
12'hf45,
12'hf84,
12'hfe2,
12'h01c,
12'h020,
12'hff7,
12'hfb4,
12'hf6c,
12'hf2a,
12'hee4,
12'he86,
12'he1a,
12'hdc5,
12'hd97,
12'hda4,
12'hdfb,
12'he7b,
12'heee,
12'hf28,
12'hf29,
12'hefe,
12'hed6,
12'hecd,
12'hed0,
12'hec4,
12'he84,
12'he3f,
12'he3c,
12'he66,
12'hea0,
12'hed5,
12'hef7,
12'hf19,
12'hf17,
12'hed7,
12'he83,
12'he65,
12'he9e,
12'hf04,
12'hf57,
12'hf69,
12'hf49,
12'hf25,
12'hf10,
12'hf1c,
12'hf4f,
12'hf8f,
12'hfaa,
12'hf92,
12'hf66,
12'hf55,
12'hf76,
12'hfbb,
12'h020,
12'h094,
12'h0e4,
12'h0df,
12'h08e,
12'h02c,
12'hfeb,
12'hfd0,
12'hfd7,
12'hfed,
12'h00f,
12'h039,
12'h05c,
12'h0b1,
12'h141,
12'h1d1,
12'h225,
12'h21d,
12'h1d8,
12'h190,
12'h159,
12'h12c,
12'h125,
12'h175,
12'h203,
12'h27a,
12'h2a6,
12'h2b4,
12'h2e8,
12'h31a,
12'h2fc,
12'h284,
12'h1ef,
12'h18e,
12'h177,
12'h1b5,
12'h22c,
12'h295,
12'h2c9,
12'h2ba,
12'h27b,
12'h221,
12'h1ba,
12'h168,
12'h131,
12'h106,
12'h0cb,
12'h083,
12'h05d,
12'h072,
12'h0b5,
12'h10a,
12'h153,
12'h168,
12'h12a,
12'h0a6,
12'h01f,
12'hfc6,
12'hf8c,
12'hf4f,
12'heef,
12'he92,
12'he74,
12'hea4,
12'hf04,
12'hf65,
12'hfc9,
12'h01b,
12'h01a,
12'hfb5,
12'hf2d,
12'hed6,
12'heb1,
12'he8e,
12'he62,
12'he4d,
12'he69,
12'head,
12'hee3,
12'hef9,
12'hf01,
12'hee8,
12'he9f,
12'he36,
12'hdf7,
12'he22,
12'he87,
12'hed8,
12'hf08,
12'hf28,
12'hf41,
12'hf47,
12'hf33,
12'hf1b,
12'hf14,
12'hf14,
12'hf0e,
12'hf0e,
12'hf27,
12'hf4a,
12'hf6d,
12'hf9f,
12'hfc4,
12'hfb9,
12'hf82,
12'hf4f,
12'hf55,
12'hf8f,
12'hfcd,
12'hfe6,
12'hfe0,
12'hfe1,
12'h017,
12'h07c,
12'h0d4,
12'h102,
12'h10d,
12'h114,
12'h111,
12'h0f9,
12'h0f4,
12'h113,
12'h143,
12'h13f,
12'h109,
12'h0df,
12'h0cf,
12'h0be,
12'h0b9,
12'h0d4,
12'h0f0,
12'h0f0,
12'h0cb,
12'h0a2,
12'h093,
12'h09a,
12'h0b1,
12'h0c0,
12'h0c5,
12'h0ab,
12'h056,
12'hff9,
12'hfd2,
12'hfe7,
12'h006,
12'h00a,
12'h010,
12'h024,
12'h01d,
12'hffd,
12'hfe5,
12'hfe1,
12'hfdd,
12'hfc3,
12'hf92,
12'hf51,
12'hf0c,
12'hece,
12'he9d,
12'he87,
12'he8b,
12'he8f,
12'heab,
12'hef8,
12'hf35,
12'hf2d,
12'heff,
12'hedb,
12'heb9,
12'he82,
12'he46,
12'he3b,
12'he7b,
12'hec5,
12'hee5,
12'hef6,
12'hf24,
12'hf64,
12'hf77,
12'hf55,
12'hf2c,
12'hf10,
12'hee2,
12'hea1,
12'he7d,
12'hea4,
12'hf05,
12'hf40,
12'hf31,
12'hf19,
12'hf43,
12'hfb2,
12'h008,
12'h02b,
12'h017,
12'hfc2,
12'hf3e,
12'hea5,
12'he43,
12'he29,
12'he47,
12'he73,
12'he84,
12'hebd,
12'hf2f,
12'hfda,
12'h093,
12'h11d,
12'h17f,
12'h1a2,
12'h186,
12'h112,
12'h040,
12'hf7b,
12'hefb,
12'hecd,
12'hef5,
12'hf60,
12'hffa,
12'h0a3,
12'h154,
12'h207,
12'h29d,
12'h301,
12'h32e,
12'h31a,
12'h29e,
12'h1bb,
12'h0b5,
12'hff3,
12'hfba,
12'h024,
12'h107,
12'h1fc,
12'h2be,
12'h331,
12'h35a,
12'h36c,
12'h371,
12'h358,
12'h304,
12'h26d,
12'h1c4,
12'h13a,
12'h0dd,
12'h0a7,
12'h0a7,
12'h0f6,
12'h165,
12'h1af,
12'h1e8,
12'h218,
12'h216,
12'h1d7,
12'h174,
12'h0f4,
12'h050,
12'hfb1,
12'hf58,
12'hf51,
12'hf7c,
12'hfa8,
12'hfc3,
12'hfc3,
12'hfa4,
12'hf71,
12'hf46,
12'hf49,
12'hf5d,
12'hf6b,
12'hf6e,
12'hf4e,
12'hf14,
12'hecf,
12'heac,
12'heb5,
12'hebc,
12'hea0,
12'he56,
12'hdfd,
12'hdbc,
12'hd9b,
12'hdae,
12'hdf4,
12'he46,
12'he77,
12'he87,
12'heaf,
12'hefe,
12'hf30,
12'hf26,
12'hf10,
12'hf1f,
12'hf48,
12'hf4b,
12'hf00,
12'he97,
12'he56,
12'he40,
12'he56,
12'hea2,
12'hf26,
12'hfc0,
12'h02d,
12'h05f,
12'h06c,
12'h072,
12'h071,
12'h043,
12'hff5,
12'hfb3,
12'hf8a,
12'hf7b,
12'hf82,
12'hfab,
12'hffd,
12'h06a,
12'h0cd,
12'h111,
12'h14e,
12'h18c,
12'h1ba,
12'h1ce,
12'h1c6,
12'h1b6,
12'h19e,
12'h17a,
12'h152,
12'h142,
12'h15b,
12'h174,
12'h16f,
12'h16a,
12'h191,
12'h1cd,
12'h1e1,
12'h1bb,
12'h163,
12'h0fc,
12'h0a9,
12'h07e,
12'h079,
12'h090,
12'h0c8,
12'h0f8,
12'h100,
12'h0ff,
12'h102,
12'h107,
12'h105,
12'h0ec,
12'h0ab,
12'h03d,
12'hfcc,
12'hf99,
12'hfbc,
12'h00a,
12'h03a,
12'h032,
12'h00f,
12'hfc7,
12'hf5c,
12'hef1,
12'he94,
12'he42,
12'hdf0,
12'hdbc,
12'hdba,
12'hddd,
12'he08,
12'he3c,
12'he86,
12'hec1,
12'heda,
12'heca,
12'he94,
12'he5c,
12'he29,
12'he0b,
12'hde6,
12'hdb6,
12'hdae,
12'hde3,
12'he4c,
12'hea4,
12'heb6,
12'he9f,
12'he95,
12'he9c,
12'he85,
12'he5e,
12'he57,
12'he65,
12'he66,
12'he5a,
12'he6a,
12'head,
12'hf00,
12'hf29,
12'hf1d,
12'hf11,
12'hf1b,
12'hf32,
12'hf51,
12'hf7e,
12'hfb1,
12'hfc3,
12'hfba,
12'hfd7,
12'h038,
12'h0a8,
12'h0d5,
12'h0b7,
12'h063,
12'hff6,
12'hf9d,
12'hf87,
12'hfc4,
12'h020,
12'h081,
12'h0d2,
12'h11e,
12'h16c,
12'h196,
12'h1a1,
12'h1a0,
12'h1a7,
12'h19c,
12'h155,
12'h109,
12'h100,
12'h15d,
12'h204,
12'h299,
12'h2fa,
12'h341,
12'h376,
12'h363,
12'h309,
12'h2a5,
12'h251,
12'h210,
12'h1f7,
12'h207,
12'h228,
12'h249,
12'h268,
12'h27b,
12'h266,
12'h22a,
12'h1d6,
12'h179,
12'h131,
12'h105,
12'h0df,
12'h0ba,
12'h0ae,
12'h0be,
12'h0da,
12'h11c,
12'h169,
12'h17a,
12'h149,
12'h0d7,
12'h03b,
12'hfa6,
12'hf39,
12'hefa,
12'heca,
12'heb0,
12'heb3,
12'hecb,
12'hf10,
12'hf62,
12'hf9b,
12'hfb8,
12'hfb1,
12'hf87,
12'hf37,
12'hee3,
12'hea5,
12'he74,
12'he47,
12'he2b,
12'he49,
12'he90,
12'hee6,
12'hf2b,
12'hf3a,
12'hf1e,
12'heda,
12'he8f,
12'he72,
12'he87,
12'heaf,
12'hed4,
12'hefc,
12'hf21,
12'hf34,
12'hf2b,
12'hf28,
12'hf49,
12'hf6f,
12'hf84,
12'hf7f,
12'hf78,
12'hf6f,
12'hf64,
12'hf7a,
12'hfa5,
12'hfcb,
12'hfe6,
12'hfe0,
12'hfd2,
12'hfd3,
12'hfdb,
12'hfe8,
12'hfe7,
12'hfe2,
12'hfff,
12'h03b,
12'h080,
12'h0af,
12'h0c9,
12'h0e7,
12'h0f6,
12'h0f2,
12'h0f9,
12'h113,
12'h132,
12'h13a,
12'h121,
12'h0f7,
12'h0c9,
12'h0ab,
12'h0aa,
12'h0c1,
12'h0cb,
12'h0bc,
12'h0a9,
12'h097,
12'h07e,
12'h071,
12'h090,
12'h0c6,
12'h0ef,
12'h0e2,
12'h099,
12'h03c,
12'hff4,
12'hfcd,
12'hfb8,
12'hfcb,
12'h011,
12'h042,
12'h045,
12'h028,
12'h009,
12'h004,
12'hff8,
12'hfdd,
12'hfb7,
12'hf6e,
12'hf06,
12'he95,
12'he56,
12'he61,
12'he83,
12'he96,
12'hea2,
12'hec5,
12'hef7,
12'hf14,
12'hf10,
12'hefb,
12'heec,
12'hed7,
12'he9d,
12'he6d,
12'he78,
12'hea0,
12'heb4,
12'heab,
12'hebb,
12'hef3,
12'hf2a,
12'hf45,
12'hf55,
12'hf7c,
12'hf93,
12'hf5a,
12'hef1,
12'hea4,
12'he9a,
12'heb5,
12'hec6,
12'hec9,
12'hee1,
12'hf2a,
12'hf8c,
12'hfea,
12'h030,
12'h048,
12'h020,
12'hf9b,
12'hef5,
12'he7d,
12'he4b,
12'he76,
12'hebe,
12'heff,
12'hf47,
12'hfa3,
12'h025,
12'h0a3,
12'h122,
12'h19c,
12'h1c8,
12'h183,
12'h0bd,
12'hfcd,
12'hf1f,
12'heda,
12'hef5,
12'hf4c,
12'hfc6,
12'h045,
12'h0c8,
12'h173,
12'h240,
12'h302,
12'h373,
12'h361,
12'h2d6,
12'h1ee,
12'h0e1,
12'h011,
12'hfcb,
12'h02f,
12'h0ff,
12'h1ca,
12'h266,
12'h2d3,
12'h328,
12'h364,
12'h36c,
12'h33c,
12'h2d5,
12'h238,
12'h192,
12'h121,
12'h0f3,
12'h0ee,
12'h0fd,
12'h125,
12'h164,
12'h19a,
12'h1cf,
12'h201,
12'h20e,
12'h1e6,
12'h18f,
12'h10e,
12'h07d,
12'h008,
12'hfcf,
12'hfd9,
12'hffc,
12'h006,
12'hff5,
12'hfc5,
12'hf80,
12'hf42,
12'hf2b,
12'hf3e,
12'hf5a,
12'hf5c,
12'hf45,
12'hf0a,
12'heb0,
12'he69,
12'he5f,
12'he95,
12'hed1,
12'hed2,
12'he94,
12'he2d,
12'hdd8,
12'hdb7,
12'hdd1,
12'he18,
12'he5b,
12'he8a,
12'he9f,
12'heb8,
12'hee2,
12'hef6,
12'hef6,
12'heee,
12'hef4,
12'hefa,
12'hedb,
12'he99,
12'he50,
12'he3c,
12'he5a,
12'he8d,
12'heda,
12'hf20,
12'hf68,
12'hfc4,
12'h026,
12'h078,
12'h09b,
12'h08e,
12'h047,
12'hfe8,
12'hfbc,
12'hfc1,
12'hfca,
12'hfd2,
12'hfea,
12'h011,
12'h034,
12'h058,
12'h098,
12'h0fb,
12'h16f,
12'h1bb,
12'h1cf,
12'h1cb,
12'h1cd,
12'h1d9,
12'h1d1,
12'h1b3,
12'h182,
12'h14c,
12'h130,
12'h12e,
12'h140,
12'h169,
12'h1b1,
12'h1e2,
12'h1c3,
12'h162,
12'h0ec,
12'h0a5,
12'h09c,
12'h0b7,
12'h0d3,
12'h0e4,
12'h0fb,
12'h104,
12'h0fd,
12'h0f4,
12'h0f9,
12'h0fe,
12'h0d5,
12'h07b,
12'h018,
12'hfd7,
12'hfbc,
12'hfc9,
12'hff1,
12'h01d,
12'h030,
12'hffc,
12'hf7f,
12'hef2,
12'he98,
12'he62,
12'he3a,
12'he28,
12'he22,
12'he1e,
12'he15,
12'he2a,
12'he6d,
12'hec3,
12'hf08,
12'hefc,
12'he97,
12'he2a,
12'hdee,
12'hdc2,
12'hda6,
12'hdaa,
12'hdd4,
12'he1d,
12'he59,
12'he82,
12'he91,
12'hea3,
12'hec4,
12'hec9,
12'heaf,
12'he69,
12'he16,
12'hddd,
12'hddc,
12'he28,
12'he97,
12'hef8,
12'hf15,
12'hede,
12'he90,
12'he7b,
12'hea3,
12'heda,
12'hf10,
12'hf2a,
12'hf36,
12'hf5a,
12'hfa8,
12'h02d,
12'h0d1,
12'h14d,
12'h152,
12'h0d5,
12'h024,
12'hf91,
12'hf3b,
12'hf2a,
12'hf59,
12'hfa7,
12'hff6,
12'h046,
12'h0b1,
12'h152,
12'h1ff,
12'h242,
12'h1fc,
12'h181,
12'h121,
12'h10a,
12'h11f,
12'h152,
12'h1ae,
12'h223,
12'h286,
12'h2a8,
12'h2c7,
12'h317,
12'h35d,
12'h362,
12'h31e,
12'h2bb,
12'h275,
12'h26e,
12'h290,
12'h2a4,
12'h2a7,
12'h27e,
12'h230,
12'h1dd,
12'h193,
12'h172,
12'h175,
12'h182,
12'h182,
12'h170,
12'h15a,
12'h13a,
12'h135,
12'h14f,
12'h162,
12'h155,
12'h108,
12'h089,
12'h01c,
12'hfe5,
12'hfce,
12'hfb4,
12'hf8d,
12'hf60,
12'hf50,
12'hf75,
12'hfae,
12'hfda,
12'hfe8,
12'hfbb,
12'hf5b,
12'hed3,
12'he51,
12'he18,
12'he25,
12'he50,
12'he52,
12'he46,
12'he66,
12'heb6,
12'hf11,
12'hf2c,
12'hf24,
12'hf03,
12'hec9,
12'he78,
12'he20,
12'he18,
12'he4d,
12'he98,
12'heca,
12'heda,
12'hf03,
12'hf22,
12'hf2b,
12'hf23,
12'hf16,
12'hf09,
12'hedf,
12'hebf,
12'hed7,
12'hf40,
12'hfc3,
12'hffd,
12'hfd2,
12'hf7b,
12'hf42,
12'hf33,
12'hf56,
12'hfa0,
12'hff7,
12'h035,
12'h038,
12'h005,
12'hfe9,
12'h01c,
12'h08a,
12'h0fd,
12'h13b,
12'h146,
12'h12f,
12'h0f8,
12'h0d8,
12'h0fc,
12'h15b,
12'h197,
12'h174,
12'h116,
12'h0b9,
12'h093,
12'h095,
12'h0c2,
12'h10f,
12'h13d,
12'h12d,
12'h0dd,
12'h083,
12'h055,
12'h064,
12'h0a2,
12'h0ce,
12'h0c8,
12'h09c,
12'h05f,
12'h033,
12'h012,
12'hffc,
12'h007,
12'h022,
12'h02e,
12'h023,
12'h003,
12'hfe3,
12'hfd7,
12'hfbe,
12'hf91,
12'hf6e,
12'hf41,
12'heee,
12'he91,
12'he5a,
12'he4d,
12'he4e,
12'he61,
12'he8e,
12'hed3,
12'hf0c,
12'hf0e,
12'hee5,
12'hea7,
12'he6c,
12'he4b,
12'he45,
12'he43,
12'he46,
12'he7e,
12'hee3,
12'hf2c,
12'hf40,
12'hf3f,
12'hf44,
12'hf39,
12'heff,
12'hec8,
12'hec6,
12'hef7,
12'hf2d,
12'hf54,
12'hf8b,
12'hfbb,
12'hfad,
12'hf59,
12'hf0a,
12'hefa,
12'hf15,
12'hf33,
12'hf3c,
12'hf47,
12'hf55,
12'hf55,
12'hf4f,
12'hf3c,
12'hf1d,
12'hef1,
12'heb4,
12'he90,
12'heae,
12'hf1c,
12'hfd8,
12'h09a,
12'h12b,
12'h18e,
12'h1c8,
12'h1d0,
12'h17f,
12'h0d5,
12'h002,
12'hf42,
12'hecc,
12'heab,
12'hf08,
12'hfcb,
12'h096,
12'h143,
12'h1cd,
12'h25c,
12'h2d1,
12'h2f5,
12'h2b7,
12'h22c,
12'h180,
12'h0ad,
12'hff3,
12'hfcd,
12'h06e,
12'h183,
12'h274,
12'h303,
12'h339,
12'h33c,
12'h32f,
12'h314,
12'h2f4,
12'h2bd,
12'h24c,
12'h1ad,
12'h113,
12'h09f,
12'h06f,
12'h0a4,
12'h130,
12'h1c7,
12'h208,
12'h1e9,
12'h19d,
12'h14f,
12'h0fe,
12'h0bf,
12'h0ae,
12'h096,
12'h058,
12'h00f,
12'hfe0,
12'hff4,
12'h033,
12'h06e,
12'h086,
12'h04b,
12'hfb1,
12'heff,
12'he85,
12'he59,
12'he81,
12'hee9,
12'hf47,
12'hf61,
12'hf35,
12'hf01,
12'heff,
12'hf1f,
12'hf28,
12'hf07,
12'hec0,
12'he4f,
12'hdda,
12'hda5,
12'hddb,
12'he67,
12'hf06,
12'hf7c,
12'hfa5,
12'hf81,
12'hf29,
12'hedc,
12'heea,
12'hf51,
12'hfb3,
12'hfc1,
12'hf73,
12'hee7,
12'he6a,
12'he39,
12'he5d,
12'hed4,
12'hf66,
12'hfe4,
12'h049,
12'h08b,
12'h09f,
12'h093,
12'h096,
12'h0a4,
12'h089,
12'h03b,
12'hfd6,
12'hf8d,
12'hf76,
12'hf87,
12'hfd8,
12'h064,
12'h0e6,
12'h12f,
12'h13c,
12'h124,
12'h116,
12'h123,
12'h154,
12'h1ab,
12'h201,
12'h216,
12'h1c8,
12'h151,
12'h100,
12'h0e8,
12'h0fd,
12'h125,
12'h149,
12'h143,
12'h0f5,
12'h079,
12'h01d,
12'h01c,
12'h071,
12'h0d1,
12'h0f9,
12'h0d1,
12'h075,
12'h037,
12'h035,
12'h05b,
12'h094,
12'h0b5,
12'h0ab,
12'h058,
12'hfbc,
12'hf34,
12'hf18,
12'hf5d,
12'hfb4,
12'hfe1,
12'hfdf,
12'hfaf,
12'hf62,
12'hf29,
12'hf27,
12'hf23,
12'hed5,
12'he37,
12'hd95,
12'hd41,
12'hd49,
12'hd9a,
12'he11,
12'he87,
12'heda,
12'hee4,
12'hebb,
12'he83,
12'he54,
12'he4a,
12'he50,
12'he45,
12'he12,
12'hdd9,
12'hde5,
12'he44,
12'hec5,
12'hf1d,
12'hf1e,
12'hef0,
12'hec5,
12'hea0,
12'he95,
12'hea8,
12'hec4,
12'hee2,
12'hef2,
12'hefe,
12'hf13,
12'hf2f,
12'hf38,
12'hf19,
12'hefb,
12'hef4,
12'hf07,
12'hf40,
12'hf7f,
12'hfa1,
12'hfa1,
12'hf9d,
12'hfd3,
12'h062,
12'h117,
12'h18b,
12'h174,
12'h0e7,
12'h02c,
12'hf87,
12'hf4c,
12'hf96,
12'h02a,
12'h09e,
12'h0c5,
12'h0d9,
12'h11c,
12'h19f,
12'h224,
12'h261,
12'h254,
12'h211,
12'h1a0,
12'h117,
12'h0ca,
12'h104,
12'h1ad,
12'h262,
12'h2c8,
12'h2e9,
12'h2f7,
12'h304,
12'h2fd,
12'h2df,
12'h2b0,
12'h25b,
12'h1eb,
12'h1a3,
12'h1a1,
12'h1db,
12'h22f,
12'h25c,
12'h24c,
12'h209,
12'h1a3,
12'h14a,
12'h123,
12'h11a,
12'h101,
12'h0bc,
12'h064,
12'h02e,
12'h039,
12'h074,
12'h0b5,
12'h0e2,
12'h0e9,
12'h0b2,
12'h03a,
12'hfa9,
12'hf31,
12'heef,
12'hecd,
12'heab,
12'he96,
12'heb6,
12'hf06,
12'hf58,
12'hf89,
12'hf98,
12'hf83,
12'hf4c,
12'hf0a,
12'hed4,
12'hebd,
12'hea7,
12'he72,
12'he35,
12'he2f,
12'he7b,
12'hedc,
12'hf09,
12'hf04,
12'heec,
12'hec7,
12'he9c,
12'he7e,
12'he95,
12'hed9,
12'hf11,
12'hf29,
12'hf31,
12'hf39,
12'hf34,
12'hf1e,
12'hf2a,
12'hf5c,
12'hf70,
12'hf48,
12'hf1f,
12'hf37,
12'hf8a,
12'hfde,
12'h000,
12'hff6,
12'hfd2,
12'hfae,
12'hf9f,
12'hfb2,
12'hfef,
12'h031,
12'h047,
12'h02c,
12'h008,
12'h015,
12'h069,
12'h0e4,
12'h142,
12'h163,
12'h150,
12'h116,
12'h0df,
12'h0e0,
12'h11f,
12'h178,
12'h1a5,
12'h17b,
12'h127,
12'h0f8,
12'h105,
12'h132,
12'h157,
12'h163,
12'h14e,
12'h11b,
12'h0d8,
12'h0a1,
12'h09f,
12'h0d8,
12'h10d,
12'h104,
12'h0cc,
12'h094,
12'h078,
12'h06f,
12'h061,
12'h04e,
12'h03d,
12'h01d,
12'hff6,
12'hfd2,
12'hfc5,
12'hfcf,
12'hfc9,
12'hfaf,
12'hf88,
12'hf56,
12'hf22,
12'heed,
12'hecb,
12'hec5,
12'hebe,
12'he94,
12'he50,
12'he2c,
12'he3b,
12'he57,
12'he62,
12'he64,
12'he77,
12'he98,
12'hea1,
12'he95,
12'he9c,
12'hebf,
12'hed5,
12'hec6,
12'heb6,
12'hebe,
12'hed5,
12'heea,
12'heed,
12'heeb,
12'hee4,
12'hebb,
12'he7c,
12'he56,
12'he69,
12'he98,
12'hea7,
12'he91,
12'he96,
12'hedf,
12'hf55,
12'hfd1,
12'h026,
12'h04e,
12'h03e,
12'hfe5,
12'hf5e,
12'hedd,
12'he80,
12'he49,
12'he33,
12'he44,
12'he9a,
12'hf44,
12'h012,
12'h0b5,
12'h10a,
12'h12c,
12'h13d,
12'h139,
12'h0fd,
12'h06b,
12'hfaf,
12'hf13,
12'hec4,
12'hece,
12'hf30,
12'hfd5,
12'h09d,
12'h178,
12'h24d,
12'h2f8,
12'h369,
12'h3a0,
12'h382,
12'h2f3,
12'h1ff,
12'h0ef,
12'h021,
12'hfe7,
12'h04f,
12'h112,
12'h1cb,
12'h24c,
12'h29a,
12'h2cc,
12'h2fb,
12'h315,
12'h30f,
12'h2ef,
12'h2a9,
12'h238,
12'h1ba,
12'h154,
12'h116,
12'h105,
12'h119,
12'h131,
12'h145,
12'h157,
12'h15a,
12'h161,
12'h18c,
12'h1c7,
12'h1ca,
12'h172,
12'h0e4,
12'h069,
12'h022,
12'hff4,
12'hfc2,
12'hf91,
12'hf63,
12'hf2c,
12'hee7,
12'heb4,
12'hebb,
12'hef5,
12'hf48,
12'hfa1,
12'hfda,
12'hfc4,
12'hf6b,
12'hf13,
12'heee,
12'heea,
12'hed2,
12'he8f,
12'he3d,
12'hdfc,
12'hdc7,
12'hda5,
12'hdc2,
12'he3e,
12'heda,
12'hf38,
12'hf44,
12'hf29,
12'hf1a,
12'hf12,
12'hf05,
12'hf06,
12'hf10,
12'hefb,
12'heb0,
12'he5e,
12'he53,
12'he92,
12'hedd,
12'hf08,
12'hf2f,
12'hf74,
12'hfc0,
12'hfe9,
12'hffd,
12'h02d,
12'h06b,
12'h061,
12'hff5,
12'hf75,
12'hf3f,
12'hf6c,
12'hfbf,
12'h00a,
12'h05c,
12'h0a8,
12'h0ca,
12'h0c5,
12'h0cc,
12'h10b,
12'h168,
12'h1a2,
12'h1b4,
12'h1a8,
12'h187,
12'h147,
12'h0f8,
12'h0da,
12'h102,
12'h138,
12'h143,
12'h145,
12'h175,
12'h1c9,
12'h1f1,
12'h1ba,
12'h153,
12'h0fa,
12'h0b7,
12'h082,
12'h064,
12'h076,
12'h0a7,
12'h0c0,
12'h0ba,
12'h0aa,
12'h0ac,
12'h0c9,
12'h0dd,
12'h0ca,
12'h08e,
12'h037,
12'hfdf,
12'hfa4,
12'hf99,
12'hfa7,
12'hfa3,
12'hf71,
12'hf1b,
12'hece,
12'hea8,
12'hea7,
12'hea7,
12'he8e,
12'he60,
12'he33,
12'he29,
12'he4a,
12'he8b,
12'hed0,
12'hef7,
12'hede,
12'he83,
12'he15,
12'hdd9,
12'hddf,
12'hdfe,
12'he08,
12'he00,
12'he13,
12'he45,
12'he8a,
12'hec1,
12'hed7,
12'hecb,
12'he9c,
12'he55,
12'he07,
12'hdd4,
12'hdc7,
12'hdc5,
12'hdce,
12'hdfc,
12'he4b,
12'he9c,
12'hecc,
12'hedd,
12'hee0,
12'hecf,
12'hea8,
12'he8f,
12'heb9,
12'hf27,
12'hf9d,
12'hfe1,
12'hff5,
12'h001,
12'h01b,
12'h034,
12'h035,
12'h019,
12'hfed,
12'hfb8,
12'hf93,
12'hf97,
12'hfd6,
12'h040,
12'h0b3,
12'h11a,
12'h168,
12'h19a,
12'h1a6,
12'h19a,
12'h193,
12'h198,
12'h190,
12'h16e,
12'h14b,
12'h15e,
12'h1bf,
12'h253,
12'h2e8,
12'h352,
12'h37d,
12'h35b,
12'h2f0,
12'h268,
12'h209,
12'h1f8,
12'h223,
12'h25b,
12'h276,
12'h26f,
12'h24d,
12'h234,
12'h245,
12'h279,
12'h297,
12'h276,
12'h227,
12'h1d5,
12'h194,
12'h15f,
12'h141,
12'h144,
12'h154,
12'h145,
12'h106,
12'h0c1,
12'h0af,
12'h0ca,
12'h0dc,
12'h0c1,
12'h08b,
12'h04d,
12'h011,
12'hfec,
12'hff6,
12'h01b,
12'h025,
12'hfe9,
12'hf7e,
12'hf2f,
12'hf07,
12'hee7,
12'hecb,
12'hecd,
12'hef4,
12'hf0d,
12'hef7,
12'hedb,
12'hef3,
12'hf40,
12'hf76,
12'hf60,
12'hf18,
12'hece,
12'he95,
12'he5e,
12'he39,
12'he45,
12'he6f,
12'he85,
12'he74,
12'he62,
12'he78,
12'heb2,
12'heef,
12'hf2c,
12'hf73,
12'hfa3,
12'hf90,
12'hf51,
12'hf34,
12'hf50,
12'hf6b,
12'hf40,
12'hee1,
12'hea5,
12'heb5,
12'heea,
12'hf25,
12'hf72,
12'hfd0,
12'h014,
12'h01b,
12'hff9,
12'hffc,
12'h03c,
12'h09b,
12'h0e1,
12'h0ec,
12'h0cc,
12'h091,
12'h04e,
12'h027,
12'h030,
12'h066,
12'h0a5,
12'h0d2,
12'h0fe,
12'h132,
12'h158,
12'h154,
12'h135,
12'h12b,
12'h138,
12'h137,
12'h10c,
12'h0d0,
12'h0ac,
12'h0a1,
12'h095,
12'h079,
12'h05a,
12'h03e,
12'h023,
12'h006,
12'hff6,
12'h00a,
12'h04f,
12'h0a2,
12'h0cd,
12'h0b9,
12'h077,
12'h038,
12'h019,
12'h00b,
12'hff9,
12'hfc9,
12'hf6a,
12'heea,
12'he73,
12'he3c,
12'he5a,
12'hea5,
12'hee9,
12'hf0d,
12'hf1a,
12'hf12,
12'hef4,
12'hec8,
12'hea4,
12'he99,
12'he9d,
12'he89,
12'he59,
12'he38,
12'he4d,
12'he8e,
12'hecd,
12'hf00,
12'hf31,
12'hf54,
12'hf48,
12'hf0a,
12'hec9,
12'heb4,
12'hec5,
12'hed7,
12'hed8,
12'hecb,
12'heae,
12'he82,
12'he6c,
12'he9a,
12'heff,
12'hf57,
12'hf77,
12'hf67,
12'hf58,
12'hf5f,
12'hf5d,
12'hf4b,
12'hf2d,
12'hf0d,
12'hee8,
12'heb4,
12'hea2,
12'heee,
12'hfa0,
12'h06d,
12'h0fe,
12'h13b,
12'h140,
12'h123,
12'h0f8,
12'h0c6,
12'h099,
12'h05c,
12'hfee,
12'hf7a,
12'hf4e,
12'hf90,
12'h016,
12'h0ad,
12'h15a,
12'h21e,
12'h2ca,
12'h31f,
12'h324,
12'h300,
12'h2bb,
12'h236,
12'h16f,
12'h0bb,
12'h077,
12'h0cc,
12'h183,
12'h236,
12'h2b5,
12'h2eb,
12'h2eb,
12'h2d5,
12'h2bf,
12'h2b4,
12'h28a,
12'h227,
12'h1b2,
12'h148,
12'h100,
12'h0ee,
12'h11e,
12'h17c,
12'h1c7,
12'h1bf,
12'h15e,
12'h0e6,
12'h0a7,
12'h0a7,
12'h0af,
12'h0a1,
12'h077,
12'h041,
12'h00e,
12'hfef,
12'h007,
12'h048,
12'h06c,
12'h03e,
12'hfbd,
12'hf1b,
12'he9d,
12'he74,
12'heb6,
12'hf42,
12'hfbd,
12'hfdd,
12'hfa4,
12'hf4f,
12'hf30,
12'hf50,
12'hf73,
12'hf66,
12'hf16,
12'hea9,
12'he36,
12'hdd3,
12'hdbe,
12'he13,
12'he99,
12'hef3,
12'hf07,
12'hefc,
12'hf02,
12'hf1c,
12'hf37,
12'hf60,
12'hf8d,
12'hf89,
12'hf3c,
12'hecc,
12'he72,
12'he3e,
12'he27,
12'he31,
12'he73,
12'hef9,
12'hf8f,
12'hff0,
12'h019,
12'h034,
12'h056,
12'h06e,
12'h06b,
12'h047,
12'h00a,
12'hfc6,
12'hf85,
12'hf64,
12'hf7d,
12'hfc2,
12'h007,
12'h02c,
12'h02a,
12'h031,
12'h06a,
12'h0cd,
12'h14a,
12'h1c5,
12'h20f,
12'h202,
12'h1a3,
12'h134,
12'h0ec,
12'h0d7,
12'h0e1,
12'h0ed,
12'h0f5,
12'h0f4,
12'h0ed,
12'h0d7,
12'h0c4,
12'h0d8,
12'h107,
12'h134,
12'h129,
12'h0e0,
12'h08f,
12'h05c,
12'h05a,
12'h078,
12'h09a,
12'h0a2,
12'h085,
12'h053,
12'h00a,
12'hfc4,
12'hf9e,
12'hf99,
12'hfb4,
12'hfdb,
12'hffc,
12'h008,
12'hfff,
12'hfeb,
12'hfc4,
12'hf84,
12'hf27,
12'hea5,
12'he22,
12'hdc2,
12'hd9b,
12'hdb3,
12'hdec,
12'he36,
12'hea7,
12'hf25,
12'hf66,
12'hf4c,
12'hf01,
12'hebd,
12'he89,
12'he42,
12'hdf1,
12'hdd6,
12'he01,
12'he3f,
12'he6d,
12'he92,
12'hec1,
12'hf08,
12'hf41,
12'hf54,
12'hf51,
12'hf46,
12'hf35,
12'hf0b,
12'hee1,
12'hedc,
12'hef3,
12'hf03,
12'hef6,
12'heda,
12'hebb,
12'he94,
12'he77,
12'he92,
12'heef,
12'hf6c,
12'hfc0,
12'hfda,
12'hfec,
12'h011,
12'h063,
12'h0b0,
12'h0c4,
12'h0a4,
12'h04b,
12'hfd3,
12'hf71,
12'hf63,
12'hfc1,
12'h049,
12'h0c3,
12'h11d,
12'h15e,
12'h18b,
12'h19c,
12'h1a3,
12'h1ae,
12'h1bb,
12'h1a6,
12'h152,
12'h0e7,
12'h0b9,
12'h106,
12'h1a0,
12'h23f,
12'h2bf,
12'h2ff,
12'h30f,
12'h2f4,
12'h2bc,
12'h292,
12'h274,
12'h26b,
12'h260,
12'h235,
12'h1f0,
12'h1a4,
12'h18e,
12'h1b9,
12'h1f2,
12'h204,
12'h1d0,
12'h187,
12'h15e,
12'h146,
12'h138,
12'h12b,
12'h113,
12'h0f1,
12'h0bd,
12'h083,
12'h04d,
12'h017,
12'hfde,
12'hf8d,
12'hf37,
12'hf06,
12'hf0c,
12'hf4b,
12'hfa8,
12'h002,
12'h036,
12'h031,
12'h008,
12'hfd6,
12'hfa0,
12'hf5c,
12'hefc,
12'he93,
12'he47,
12'he33,
12'he47,
12'he6f,
12'hea8,
12'hee9,
12'hf22,
12'hf33,
12'hf29,
12'hf22,
12'hf21,
12'hf2e,
12'hf2c,
12'hf0e,
12'hee8,
12'hec7,
12'heb9,
12'heba,
12'hedd,
12'hf1f,
12'hf51,
12'hf42,
12'hefc,
12'hec5,
12'hed6,
12'hf22,
12'hf6f,
12'hfa0,
12'hfa1,
12'hf6a,
12'hf2b,
12'hf18,
12'hf4f,
12'hfb8,
12'h006,
12'h016,
12'hff3,
12'hfc1,
12'hf9d,
12'hf95,
12'hfbb,
12'h00e,
12'h06b,
12'h0a2,
12'h0b3,
12'h0b5,
12'h0ca,
12'h0fc,
12'h12b,
12'h12b,
12'h0fe,
12'h0d4,
12'h0b9,
12'h0aa,
12'h0b3,
12'h0e0,
12'h11b,
12'h13f,
12'h13c,
12'h11c,
12'h107,
12'h0f7,
12'h0d1,
12'h094,
12'h047,
12'h023,
12'h02f,
12'h03c,
12'h040,
12'h049,
12'h065,
12'h08c,
12'h0aa,
12'h0b8,
12'h0c2,
12'h0c4,
12'h0a4,
12'h060,
12'h01a,
12'hfdd,
12'hfb5,
12'hfa6,
12'hf95,
12'hf7d,
12'hf4c,
12'hf0d,
12'hedb,
12'hed7,
12'hf0e,
12'hf4c,
12'hf5b,
12'hf3e,
12'hf1b,
12'hefe,
12'hee0,
12'hec5,
12'hebc,
12'hebe,
12'hea9,
12'he7e,
12'he53,
12'he65,
12'heaf,
12'hef8,
12'hf42,
12'hf6a,
12'hf71,
12'hf4d,
12'hf03,
12'hee5,
12'hf04,
12'hf35,
12'hf3b,
12'hf0f,
12'heee,
12'hef6,
12'hf0f,
12'hf16,
12'hf0f,
12'hf11,
12'hefa,
12'head,
12'he6c,
12'he85,
12'hef2,
12'hf60,
12'hf7b,
12'hf51,
12'hf1a,
12'hef1,
12'hee2,
12'heff,
12'hf3c,
12'hf72,
12'hf86,
12'hf8e,
12'hfb6,
12'h003,
12'h063,
12'h0ad,
12'h0c3,
12'h092,
12'h02d,
12'hfc5,
12'hf80,
12'hf88,
12'hfc7,
12'h01c,
12'h074,
12'h0be,
12'h108,
12'h15e,
12'h1c3,
12'h231,
12'h28a,
12'h293,
12'h23b,
12'h1a9,
12'h117,
12'h0ce,
12'h0ef,
12'h16c,
12'h207,
12'h28b,
12'h2db,
12'h2e1,
12'h2c4,
12'h2a8,
12'h296,
12'h28a,
12'h267,
12'h223,
12'h1ce,
12'h189,
12'h173,
12'h188,
12'h1a9,
12'h1ac,
12'h183,
12'h147,
12'h10b,
12'h0f9,
12'h110,
12'h122,
12'h11f,
12'h0f3,
12'h0a1,
12'h04c,
12'h01e,
12'h037,
12'h06f,
12'h086,
12'h059,
12'hfe6,
12'hf5b,
12'heea,
12'hea5,
12'hea6,
12'heea,
12'hf5b,
12'hfbd,
12'hfc3,
12'hf7e,
12'hf35,
12'hf28,
12'hf45,
12'hf4b,
12'hf2b,
12'hedb,
12'he65,
12'hdea,
12'hd9d,
12'hdb4,
12'he22,
12'heac,
12'hf0f,
12'hf24,
12'hf06,
12'heef,
12'heec,
12'hf00,
12'hf1f,
12'hf29,
12'hf11,
12'hecc,
12'he7c,
12'he63,
12'he8c,
12'heeb,
12'hf5a,
12'hfb6,
12'hfe4,
12'hfe1,
12'hfcc,
12'hfd2,
12'h019,
12'h06f,
12'h077,
12'h027,
12'hfc1,
12'hf80,
12'hf76,
12'hfa6,
12'hffd,
12'h047,
12'h061,
12'h044,
12'h01a,
12'h01f,
12'h06c,
12'h0ef,
12'h16f,
12'h1ac,
12'h198,
12'h157,
12'h119,
12'h106,
12'h11d,
12'h142,
12'h153,
12'h134,
12'h0fe,
12'h0da,
12'h0d3,
12'h0e2,
12'h0e8,
12'h0e0,
12'h0d3,
12'h0af,
12'h087,
12'h075,
12'h087,
12'h0b3,
12'h0cc,
12'h0c4,
12'h098,
12'h060,
12'h034,
12'h014,
12'h018,
12'h027,
12'h01d,
12'hfeb,
12'hf95,
12'hf54,
12'hf55,
12'hf91,
12'hfdd,
12'hffa,
12'hfcc,
12'hf60,
12'hed4,
12'he65,
12'he2d,
12'he1e,
12'he1c,
12'he13,
12'he0d,
12'he08,
12'he0e,
12'he42,
12'he8e,
12'hecb,
12'hed1,
12'hea1,
12'he7d,
12'he6d,
12'he4b,
12'he17,
12'hdf0,
12'he01,
12'he45,
12'he86,
12'heb2,
12'hef3,
12'hf59,
12'hfa3,
12'hf91,
12'hf41,
12'hf01,
12'hef1,
12'hede,
12'heb0,
12'he8d,
12'he84,
12'he9d,
12'hed5,
12'hf1a,
12'hf4c,
12'hf56,
12'hf4b,
12'hf36,
12'hf3b,
12'hf86,
12'hffc,
12'h068,
12'h09f,
12'h09f,
12'h09b,
12'h0ab,
12'h0b4,
12'h09b,
12'h046,
12'hfd7,
12'hf88,
12'hf75,
12'hfbc,
12'h056,
12'h102,
12'h196,
12'h208,
12'h244,
12'h236,
12'h1e6,
12'h17e,
12'h135,
12'h104,
12'h0d5,
12'h0b4,
12'h0cf,
12'h156,
12'h21d,
12'h2cd,
12'h336,
12'h36e,
12'h399,
12'h392,
12'h33b,
12'h2b9,
12'h23f,
12'h1ee,
12'h1c0,
12'h1ad,
12'h1b1,
12'h1b4,
12'h1bc,
12'h1df,
12'h214,
12'h246,
12'h257,
12'h247,
12'h21c,
12'h1c5,
12'h14f,
12'h0cf,
12'h068,
12'h035,
12'h03e,
12'h06d,
12'h094,
12'h09e,
12'h085,
12'h060,
12'h04e,
12'h039,
12'h00d,
12'hfd6,
12'hf9b,
12'hf63,
12'hf33,
12'hf1f,
12'hf3b,
12'hf65,
12'hf71,
12'hf3b,
12'hecb,
12'he5e,
12'he23,
12'he38,
12'he7d,
12'heb0,
12'heb1,
12'he95,
12'he7e,
12'he65,
12'he5e,
12'he83,
12'heb8,
12'hecd,
12'he97,
12'he3b,
12'he0c,
12'he24,
12'he73,
12'hed8,
12'hf17,
12'hf1d,
12'hee7,
12'he94,
12'he66,
12'he72,
12'hebb,
12'hf18,
12'hf58,
12'hf75,
12'hf71,
12'hf7b,
12'hfaf,
12'hfdf,
12'hfed,
12'hfdc,
12'hfa3,
12'hf4b,
12'hf14,
12'hf21,
12'hf66,
12'hfbd,
12'h000,
12'h041,
12'h085,
12'h0b4,
12'h0c5,
12'h0c7,
12'h0e3,
12'h114,
12'h121,
12'h0fb,
12'h0bf,
12'h0a1,
12'h0ba,
12'h0e9,
12'h10f,
12'h132,
12'h14a,
12'h149,
12'h139,
12'h11f,
12'h113,
12'h115,
12'h0f8,
12'h0b5,
12'h065,
12'h03e,
12'h053,
12'h08d,
12'h0be,
12'h0d3,
12'h0dc,
12'h0d7,
12'h0cc,
12'h0ae,
12'h085,
12'h05e,
12'h038,
12'h01c,
12'h00d,
12'h020,
12'h040,
12'h04b,
12'h043,
12'h029,
12'hffd,
12'hfa9,
12'hf38,
12'hece,
12'he8e,
12'he90,
12'hebf,
12'hf06,
12'hf54,
12'hf94,
12'hf92,
12'hf4d,
12'hf0e,
12'hef5,
12'hed9,
12'he90,
12'he39,
12'he18,
12'he43,
12'he82,
12'heb2,
12'hee1,
12'hf11,
12'hf2e,
12'hf1d,
12'hf18,
12'hf58,
12'hf9e,
12'hfaf,
12'hf80,
12'hf36,
12'hf03,
12'hed8,
12'hea3,
12'he76,
12'he60,
12'he55,
12'he41,
12'he4b,
12'heb8,
12'hf6c,
12'hffe,
12'h013,
12'hfb2,
12'hf2c,
12'heb5,
12'he66,
12'he59,
12'he8f,
12'hedf,
12'hf13,
12'hf34,
12'hf72,
12'hfef,
12'h09b,
12'h130,
12'h173,
12'h131,
12'h084,
12'hfc2,
12'hf3e,
12'hf2c,
12'hf60,
12'hfba,
12'h029,
12'h092,
12'h0f0,
12'h155,
12'h1dc,
12'h269,
12'h2b5,
12'h29c,
12'h224,
12'h190,
12'h128,
12'h111,
12'h13f,
12'h197,
12'h20f,
12'h279,
12'h2b3,
12'h2c6,
12'h2d9,
12'h2f6,
12'h305,
12'h2f1,
12'h2bb,
12'h268,
12'h202,
12'h1ae,
12'h181,
12'h171,
12'h161,
12'h140,
12'h12a,
12'h13d,
12'h171,
12'h18d,
12'h16b,
12'h13c,
12'h113,
12'h0db,
12'h088,
12'h03d,
12'h022,
12'h028,
12'h03a,
12'h03f,
12'h02d,
12'h00b,
12'hfd9,
12'hf83,
12'hf0d,
12'he90,
12'he47,
12'he71,
12'hf00,
12'hf8c,
12'hfb6,
12'hf8e,
12'hf58,
12'hf26,
12'hef5,
12'hec2,
12'hea0,
12'he89,
12'he56,
12'he13,
12'hde4,
12'hdfc,
12'he58,
12'heba,
12'hef0,
12'heef,
12'hecc,
12'he94,
12'he6e,
12'he94,
12'hf10,
12'hf93,
12'hfb6,
12'hf6c,
12'hee0,
12'he62,
12'he3b,
12'he67,
12'hee5,
12'hf7a,
12'hfd0,
12'hfcc,
12'hfa9,
12'hfbf,
12'h014,
12'h063,
12'h062,
12'h019,
12'hfb3,
12'hf71,
12'hf7e,
12'hfcb,
12'h052,
12'h0d8,
12'h109,
12'h0ce,
12'h05d,
12'h028,
12'h05c,
12'h0c8,
12'h126,
12'h155,
12'h168,
12'h176,
12'h184,
12'h17e,
12'h16f,
12'h15b,
12'h148,
12'h129,
12'h0fc,
12'h0ed,
12'h100,
12'h115,
12'h110,
12'h0f0,
12'h0d7,
12'h0cf,
12'h0d0,
12'h0ce,
12'h0cf,
12'h0d7,
12'h0c6,
12'h08e,
12'h055,
12'h047,
12'h05c,
12'h06d,
12'h05a,
12'h02a,
12'hff5,
12'hfb4,
12'hf82,
12'hf8a,
12'hfda,
12'h02c,
12'h033,
12'hff5,
12'hf93,
12'hf3b,
12'heed,
12'he92,
12'he42,
12'he02,
12'hdd3,
12'hdb8,
12'hdc6,
12'he06,
12'he68,
12'hed9,
12'hf21,
12'hf22,
12'hedf,
12'he7e,
12'he3e,
12'he2f,
12'he35,
12'he3d,
12'he3a,
12'he4c,
12'he94,
12'heea,
12'hf2d,
12'hf58,
12'hf6b,
12'hf57,
12'hef9,
12'he8f,
12'he66,
12'he83,
12'heb8,
12'hec7,
12'hece,
12'heee,
12'hf2d,
12'hf5a,
12'hf52,
12'hf46,
12'hf29,
12'hf03,
12'hefb,
12'hf27,
12'hf83,
12'hfd4,
12'hffd,
12'h00a,
12'h032,
12'h081,
12'h0cc,
12'h0d1,
12'h075,
12'hff7,
12'hf78,
12'hf33,
12'hf51,
12'hfbe,
12'h04a,
12'h0bb,
12'h10f,
12'h150,
12'h18a,
12'h1c1,
12'h1f5,
12'h21d,
12'h20d,
12'h1b8,
12'h127,
12'h0aa,
12'h097,
12'h0f3,
12'h19f,
12'h258,
12'h2ef,
12'h358,
12'h389,
12'h385,
12'h35c,
12'h311,
12'h2a3,
12'h240,
12'h1f0,
12'h1a4,
12'h164,
12'h145,
12'h16b,
12'h1c9,
12'h216,
12'h224,
12'h1f8,
12'h1be,
12'h19a,
12'h187,
12'h17b,
12'h15b,
12'h109,
12'h0a7,
12'h069,
12'h05f,
12'h077,
12'h093,
12'h08a,
12'h033,
12'hfba,
12'hf5e,
12'hf52,
12'hf93,
12'hfd1,
12'hfd8,
12'hfa4,
12'hf5d,
12'hf22,
12'hef7,
12'hef2,
12'hf05,
12'hefd,
12'hec9,
12'he88,
12'he66,
12'he6c,
12'he8e,
12'heb7,
12'hece,
12'hecf,
12'heb4,
12'he83,
12'he68,
12'he70,
12'he90,
12'heb9,
12'hec4,
12'heb6,
12'he9e,
12'he86,
12'he8c,
12'heae,
12'hed7,
12'hee8,
12'hec2,
12'hea8,
12'hecc,
12'hf2b,
12'hfb1,
12'h011,
12'h021,
12'hfec,
12'hfa2,
12'hf71,
12'hf67,
12'hf83,
12'hf97,
12'hf9a,
12'hf95,
12'hf91,
12'hfa1,
12'hfc0,
12'hff9,
12'h03a,
12'h067,
12'h07c,
12'h076,
12'h07a,
12'h09f,
12'h0f0,
12'h14e,
12'h18b,
12'h195,
12'h167,
12'h126,
12'h0ef,
12'h0d2,
12'h0ce,
12'h0da,
12'h0fd,
12'h121,
12'h136,
12'h13e,
12'h135,
12'h11e,
12'h0ef,
12'h09f,
12'h05b,
12'h050,
12'h084,
12'h0d7,
12'h107,
12'h0f9,
12'h0d3,
12'h0a8,
12'h078,
12'h04f,
12'h043,
12'h04c,
12'h056,
12'h044,
12'h015,
12'hff9,
12'h003,
12'h025,
12'h02d,
12'h008,
12'hfb9,
12'hf4b,
12'hee4,
12'heb3,
12'hec2,
12'hee5,
12'heeb,
12'hede,
12'hed3,
12'hec4,
12'hebb,
12'heca,
12'hee3,
12'heed,
12'hed1,
12'he94,
12'he6d,
12'he6b,
12'he73,
12'he88,
12'heb5,
12'hede,
12'hee8,
12'hec7,
12'heb4,
12'heee,
12'hf4d,
12'hf7f,
12'hf5c,
12'hf15,
12'heeb,
12'hed8,
12'heb3,
12'he76,
12'he41,
12'he35,
12'he6b,
12'hedc,
12'hf68,
12'hff7,
12'h04c,
12'h03b,
12'hfc7,
12'hf2e,
12'hecb,
12'heb9,
12'hed3,
12'hedc,
12'hed5,
12'hee8,
12'hf2c,
12'hfa5,
12'h049,
12'h0f3,
12'h15a,
12'h141,
12'h0b9,
12'h016,
12'hfb3,
12'hf95,
12'hfa7,
12'hfdb,
12'h012,
12'h04c,
12'h097,
12'h0fd,
12'h17a,
12'h1ff,
12'h26e,
12'h2a9,
12'h29f,
12'h246,
12'h1b2,
12'h13d,
12'h124,
12'h157,
12'h1a3,
12'h1d8,
12'h213,
12'h263,
12'h2a9,
12'h2d0,
12'h2d7,
12'h2d7,
12'h2c5,
12'h299,
12'h265,
12'h22f,
12'h20b,
12'h1df,
12'h19b,
12'h160,
12'h12b,
12'h100,
12'h0f5,
12'h112,
12'h13d,
12'h14e,
12'h134,
12'h0f4,
12'h09e,
12'h058,
12'h040,
12'h059,
12'h078,
12'h085,
12'h076,
12'h042,
12'h007,
12'hfba,
12'hf39,
12'heab,
12'he4a,
12'he37,
12'he7a,
12'hee3,
12'hf4a,
12'hfa0,
12'hfc8,
12'hfae,
12'hf6b,
12'hf30,
12'hefd,
12'hebd,
12'he71,
12'he23,
12'hdef,
12'hdff,
12'he51,
12'heb6,
12'hefe,
12'hf12,
12'hef9,
12'hebe,
12'he7f,
12'he75,
12'hec1,
12'hf41,
12'hfab,
12'hfcc,
12'hf94,
12'hf1e,
12'hec2,
12'heb3,
12'hef1,
12'hf3e,
12'hf61,
12'hf70,
12'hf89,
12'hfab,
12'hfec,
12'h04d,
12'h08c,
12'h070,
12'h017,
12'hfaa,
12'hf50,
12'hf39,
12'hf93,
12'h043,
12'h0cd,
12'h0e9,
12'h0aa,
12'h05b,
12'h041,
12'h065,
12'h0bc,
12'h119,
12'h149,
12'h144,
12'h12a,
12'h119,
12'h120,
12'h133,
12'h13a,
12'h125,
12'h103,
12'h0ed,
12'h0eb,
12'h0f5,
12'h102,
12'h104,
12'h0e7,
12'h0ba,
12'h0b3,
12'h0d7,
12'h103,
12'h116,
12'h105,
12'h0ce,
12'h079,
12'h036,
12'h027,
12'h039,
12'h042,
12'h036,
12'h015,
12'hfd4,
12'hf89,
12'hf5a,
12'hf6d,
12'hfc2,
12'h012,
12'h029,
12'hffc,
12'hfa6,
12'hf55,
12'hf11,
12'hecf,
12'he89,
12'he46,
12'he01,
12'hdc8,
12'hdd3,
12'he20,
12'he7f,
12'hec2,
12'hed6,
12'hec3,
12'he99,
12'he61,
12'he2d,
12'he2e,
12'he67,
12'he9a,
12'he9c,
12'he8d,
12'heb0,
12'hefe,
12'hf42,
12'hf66,
12'hf57,
12'hf1f,
12'hed4,
12'he87,
12'he5d,
12'he7a,
12'hedd,
12'hf2c,
12'hf23,
12'hef4,
12'hef5,
12'hf4c,
12'hfad,
12'hfc2,
12'hf94,
12'hf35,
12'hed0,
12'he8a,
12'he90,
12'hf06,
12'hfa2,
12'hff8,
12'h002,
12'h018,
12'h077,
12'h0f4,
12'h12b,
12'h0fd,
12'h08b,
12'hff9,
12'hf67,
12'hf24,
12'hf56,
12'hfd5,
12'h045,
12'h088,
12'h0d2,
12'h144,
12'h1bb,
12'h210,
12'h238,
12'h230,
12'h1ef,
12'h163,
12'h0d1,
12'h0a5,
12'h0fa,
12'h19c,
12'h231,
12'h295,
12'h2e6,
12'h331,
12'h35a,
12'h35c,
12'h33f,
12'h2f9,
12'h28d,
12'h213,
12'h1af,
12'h172,
12'h162,
12'h185,
12'h1bc,
12'h1e4,
12'h1d4,
12'h18f,
12'h15a,
12'h15b,
12'h183,
12'h192,
12'h17d,
12'h14c,
12'h0fb,
12'h0b0,
12'h07d,
12'h074,
12'h08c,
12'h085,
12'h049,
12'hfd9,
12'hf69,
12'hf48,
12'hf73,
12'hfac,
12'hfb5,
12'hf91,
12'hf48,
12'hee4,
12'he93,
12'he84,
12'hebd,
12'hf0c,
12'hf35,
12'hf28,
12'hf01,
12'hede,
12'heb8,
12'hea1,
12'hea1,
12'hea2,
12'hea1,
12'he87,
12'he60,
12'he5e,
12'he87,
12'hec0,
12'hee3,
12'hef4,
12'hf11,
12'hf1f,
12'hf0c,
12'heed,
12'heeb,
12'hefc,
12'hef4,
12'hed9,
12'hec7,
12'hed2,
12'hefa,
12'hf42,
12'hf9c,
12'hfe0,
12'hff9,
12'hfe4,
12'hfb4,
12'hf94,
12'hf90,
12'hfa0,
12'hfc3,
12'hfe7,
12'hfe9,
12'hfd7,
12'hfcd,
12'hfdb,
12'h008,
12'h042,
12'h079,
12'h09c,
12'h0ac,
12'h0b9,
12'h0c3,
12'h0d7,
12'h10a,
12'h13b,
12'h149,
12'h130,
12'h0f4,
12'h0a4,
12'h067,
12'h067,
12'h0be,
12'h133,
12'h179,
12'h173,
12'h125,
12'h0bd,
12'h05f,
12'h02d,
12'h039,
12'h083,
12'h0ca,
12'h0d3,
12'h0ab,
12'h081,
12'h083,
12'h098,
12'h098,
12'h07f,
12'h054,
12'h019,
12'hfe2,
12'hfca,
12'hfe8,
12'h02d,
12'h05a,
12'h03a,
12'hfe4,
12'hf7d,
12'hf0f,
12'heb2,
12'he85,
12'he94,
12'heb9,
12'heca,
12'hec4,
12'heaf,
12'hea4,
12'heb5,
12'hecb,
12'hed4,
12'hed9,
12'hecd,
12'heac,
12'he92,
12'he83,
12'he84,
12'he92,
12'heb7,
12'hef0,
12'hf09,
12'hf03,
12'hf10,
12'hf32,
12'hf3a,
12'hf18,
12'hef1,
12'hee4,
12'hedf,
12'heb3,
12'he6a,
12'he30,
12'he24,
12'he53,
12'hec1,
12'hf41,
12'hfb5,
12'hffe,
12'h00a,
12'hffa,
12'hfda,
12'hfa9,
12'hf56,
12'hefa,
12'heb9,
12'head,
12'heeb,
12'hf49,
12'hfc0,
12'h049,
12'h0b2,
12'h0df,
12'h0db,
12'h0c8,
12'h090,
12'h02d,
12'hfc0,
12'hf6d,
12'hf63,
12'hf9d,
12'hffa,
12'h07d,
12'h12b,
12'h1d5,
12'h231,
12'h247,
12'h255,
12'h27a,
12'h28d,
12'h24b,
12'h1d3,
12'h179,
12'h169,
12'h197,
12'h1e4,
12'h24e,
12'h2a5,
12'h2af,
12'h27f,
12'h246,
12'h23e,
12'h259,
12'h27a,
12'h299,
12'h28c,
12'h23f,
12'h1cd,
12'h178,
12'h16f,
12'h18e,
12'h18d,
12'h156,
12'h111,
12'h100,
12'h110,
12'h10e,
12'h104,
12'h0ff,
12'h0e6,
12'h0a2,
12'h05a,
12'h035,
12'h037,
12'h052,
12'h064,
12'h057,
12'hffa,
12'hf41,
12'he68,
12'hdd3,
12'hdd2,
12'he50,
12'heef,
12'hf66,
12'hfad,
12'hfc9,
12'hfc2,
12'hf9f,
12'hf68,
12'hf35,
12'hef1,
12'he81,
12'hdfa,
12'hd9e,
12'hdac,
12'he0e,
12'he75,
12'hec8,
12'hefb,
12'hf01,
12'hed6,
12'he86,
12'he55,
12'he5f,
12'heab,
12'hf12,
12'hf5e,
12'hf76,
12'hf4d,
12'hf10,
12'hedb,
12'hecf,
12'hee9,
12'hf0c,
12'hf3c,
12'hf77,
12'hfac,
12'hfd8,
12'h006,
12'h037,
12'h04e,
12'h025,
12'hfd1,
12'hf69,
12'hf2e,
12'hf57,
12'hfc9,
12'h045,
12'h096,
12'h0bb,
12'h0b7,
12'h092,
12'h06b,
12'h064,
12'h09f,
12'h11a,
12'h193,
12'h1c2,
12'h19c,
12'h14d,
12'h10d,
12'h0ef,
12'h0ec,
12'h0fa,
12'h107,
12'h102,
12'h0e1,
12'h0b2,
12'h095,
12'h0ad,
12'h0ee,
12'h130,
12'h154,
12'h130,
12'h0df,
12'h0a0,
12'h092,
12'h09d,
12'h09b,
12'h08a,
12'h074,
12'h050,
12'h023,
12'h014,
12'h01c,
12'h018,
12'hfec,
12'hfaa,
12'hf8a,
12'hf95,
12'hfac,
12'hfb6,
12'hfb4,
12'hf9f,
12'hf4b,
12'hed1,
12'he6b,
12'he31,
12'he2e,
12'he44,
12'he67,
12'he95,
12'hebd,
12'hee6,
12'hf02,
12'hf03,
12'hee0,
12'he8f,
12'he36,
12'hdfc,
12'hdf4,
12'he1c,
12'he53,
12'hea0,
12'hf19,
12'hf8b,
12'hfbd,
12'hfb7,
12'hf95,
12'hf6b,
12'hf30,
12'hedc,
12'he87,
12'he5f,
12'he80,
12'hebd,
12'hee2,
12'heeb,
12'hf09,
12'hf5d,
12'hfa0,
12'hf9b,
12'hf69,
12'hf30,
12'hf00,
12'hed9,
12'hecc,
12'hef8,
12'hf48,
12'hf7d,
12'hf89,
12'hfad,
12'h025,
12'h0a9,
12'h0dd,
12'h0bc,
12'h06e,
12'h015,
12'hfbb,
12'hf92,
12'hfb7,
12'h004,
12'h041,
12'h065,
12'h0a2,
12'h10c,
12'h17f,
12'h1db,
12'h20d,
12'h215,
12'h1d1,
12'h13e,
12'h0b8,
12'h09e,
12'h106,
12'h1a1,
12'h221,
12'h281,
12'h2e4,
12'h34e,
12'h38d,
12'h391,
12'h36c,
12'h31b,
12'h29c,
12'h206,
12'h193,
12'h166,
12'h180,
12'h1bb,
12'h1f1,
12'h204,
12'h1d8,
12'h191,
12'h15c,
12'h154,
12'h166,
12'h161,
12'h139,
12'h0f9,
12'h0ab,
12'h05f,
12'h031,
12'h02f,
12'h049,
12'h062,
12'h055,
12'h00b,
12'hfae,
12'hf77,
12'hf83,
12'hfae,
12'hfb7,
12'hf88,
12'hf30,
12'hec9,
12'he8b,
12'he8a,
12'hebb,
12'heff,
12'hf29,
12'hf20,
12'hef4,
12'hecb,
12'heab,
12'he9d,
12'hea6,
12'heab,
12'he9c,
12'he6e,
12'he45,
12'he54,
12'he8d,
12'hed0,
12'hefa,
12'hf0f,
12'hf24,
12'hf28,
12'hf0c,
12'hee5,
12'hee0,
12'hefa,
12'hf01,
12'hef1,
12'hee1,
12'hef1,
12'hf25,
12'hf67,
12'hfa7,
12'hfe2,
12'h011,
12'h00a,
12'hfc3,
12'hf62,
12'hf26,
12'hf37,
12'hf80,
12'hfd1,
12'h010,
12'h02b,
12'h026,
12'h021,
12'h038,
12'h06b,
12'h0a2,
12'h0cc,
12'h0c7,
12'h09c,
12'h074,
12'h078,
12'h0bb,
12'h115,
12'h15e,
12'h178,
12'h145,
12'h0e5,
12'h08f,
12'h07f,
12'h0c5,
12'h121,
12'h151,
12'h13f,
12'h102,
12'h0ad,
12'h052,
12'h023,
12'h04f,
12'h0bf,
12'h10e,
12'h0fe,
12'h0b7,
12'h07d,
12'h071,
12'h074,
12'h074,
12'h071,
12'h055,
12'h016,
12'hfcb,
12'hfa1,
12'hfb3,
12'hff3,
12'h02b,
12'h033,
12'hff2,
12'hf76,
12'hef9,
12'hea2,
12'he95,
12'hec6,
12'heef,
12'hede,
12'hea7,
12'he71,
12'he59,
12'he74,
12'heaa,
12'hede,
12'hefb,
12'hef1,
12'hed5,
12'hec4,
12'hebd,
12'hec0,
12'hebe,
12'hebe,
12'hecc,
12'hed5,
12'heec,
12'hf1d,
12'hf56,
12'hf62,
12'hf32,
12'hef4,
12'hed6,
12'hec8,
12'hea5,
12'he74,
12'he53,
12'he69,
12'heb7,
12'hf1b,
12'hf88,
12'hff6,
12'h03c,
12'h03b,
12'h000,
12'hfb5,
12'hf65,
12'hf03,
12'heb8,
12'hea6,
12'hecd,
12'hf1a,
12'hf76,
12'hfe8,
12'h054,
12'h09e,
12'h0c4,
12'h0d2,
12'h0c1,
12'h06e,
12'hfee,
12'hf84,
12'hf68,
12'hf97,
12'hfef,
12'h05a,
12'h0e3,
12'h170,
12'h1c4,
12'h1da,
12'h1ef,
12'h239,
12'h289,
12'h27e,
12'h212,
12'h1a0,
12'h16c,
12'h184,
12'h1d1,
12'h241,
12'h2bf,
12'h2f6,
12'h2c0,
12'h250,
12'h1fe,
12'h1f9,
12'h21c,
12'h24b,
12'h27b,
12'h273,
12'h220,
12'h1c2,
12'h194,
12'h1a4,
12'h1ac,
12'h17d,
12'h132,
12'h0f7,
12'h0da,
12'h0bd,
12'h0ab,
12'h0bc,
12'h0d4,
12'h0c5,
12'h079,
12'h02d,
12'h013,
12'h021,
12'h03a,
12'h039,
12'h00b,
12'hfa4,
12'hef9,
12'he45,
12'hde2,
12'hdfb,
12'he6e,
12'hef4,
12'hf72,
12'hfc9,
12'hfd2,
12'hf93,
12'hf4e,
12'hf36,
12'hf29,
12'hef5,
12'he84,
12'he18,
12'hdfa,
12'he1f,
12'he64,
12'heb5,
12'hf0f,
12'hf4b,
12'hf3b,
12'heea,
12'he8f,
12'he5d,
12'he71,
12'hec6,
12'hf35,
12'hf90,
12'hfac,
12'hf7d,
12'hf2d,
12'hef4,
12'heeb,
12'hf12,
12'hf50,
12'hf96,
12'hfc7,
12'hfc1,
12'hfb2,
12'hfcd,
12'h001,
12'h027,
12'h011,
12'hfbd,
12'hf66,
12'hf4f,
12'hf8e,
12'h000,
12'h071,
12'h0b6,
12'h0c4,
12'h0ab,
12'h07b,
12'h05a,
12'h06d,
12'h0d1,
12'h158,
12'h1aa,
12'h19f,
12'h150,
12'h0fe,
12'h0cc,
12'h0c9,
12'h0e4,
12'h104,
12'h117,
12'h10a,
12'h0e3,
12'h0be,
12'h0c2,
12'h0ee,
12'h119,
12'h12c,
12'h121,
12'h0fb,
12'h0d4,
12'h0b5,
12'h098,
12'h06f,
12'h03b,
12'h018,
12'h004,
12'hff4,
12'hfef,
12'hfec,
12'hfe0,
12'hfcb,
12'hfbc,
12'hfb4,
12'hfaa,
12'hf96,
12'hf7a,
12'hf6b,
12'hf63,
12'hf48,
12'hf07,
12'heac,
12'he68,
12'he35,
12'he10,
12'he1c,
12'he56,
12'he96,
12'hebf,
12'hed4,
12'hed6,
12'hec0,
12'he97,
12'he4d,
12'hdff,
12'hde4,
12'he06,
12'he44,
12'he83,
12'hee9,
12'hf6d,
12'hfcf,
12'hfe4,
12'hfaf,
12'hf69,
12'hf29,
12'hed3,
12'he73,
12'he2e,
12'he32,
12'he7b,
12'hebe,
12'hef2,
12'hf3d,
12'hfa6,
12'hff0,
12'hfce,
12'hf6e,
12'hf1c,
12'heeb,
12'hed7,
12'hee1,
12'hf17,
12'hf55,
12'hf77,
12'hf85,
12'hfa0,
12'hff9,
12'h074,
12'h0c3,
12'h0c5,
12'h087,
12'h02d,
12'hfd7,
12'hfb1,
12'hfcd,
12'hffd,
12'h024,
12'h034,
12'h04c,
12'h0a2,
12'h13e,
12'h1de,
12'h236,
12'h23b,
12'h1ec,
12'h165,
12'h0f5,
12'h0cd,
12'h10a,
12'h192,
12'h20f,
12'h254,
12'h285,
12'h2db,
12'h342,
12'h389,
12'h39d,
12'h36b,
12'h2e6,
12'h241,
12'h1c4,
12'h196,
12'h1ba,
12'h206,
12'h236,
12'h224,
12'h1dd,
12'h187,
12'h153,
12'h14a,
12'h157,
12'h162,
12'h14f,
12'h119,
12'h0d4,
12'h09e,
12'h08a,
12'h08c,
12'h077,
12'h046,
12'h021,
12'h007,
12'hfdb,
12'hf9e,
12'hf85,
12'hf91,
12'hf89,
12'hf5a,
12'hf24,
12'hf06,
12'hed8,
12'he94,
12'he74,
12'he9a,
12'heea,
12'hf25,
12'hf2f,
12'hf19,
12'heef,
12'head,
12'he70,
12'he69,
12'he95,
12'heb9,
12'hea7,
12'he7d,
12'he67,
12'he74,
12'he9a,
12'hed5,
12'hf27,
12'hf6a,
12'hf71,
12'hf38,
12'hf00,
12'hefe,
12'hf1c,
12'hf3a,
12'hf45,
12'hf49,
12'hf43,
12'hf36,
12'hf45,
12'hf90,
12'h00b,
12'h064,
12'h04a,
12'hfd2,
12'hf53,
12'hf19,
12'hf38,
12'hf91,
12'hff8,
12'h040,
12'h049,
12'h029,
12'h00b,
12'h01f,
12'h06c,
12'h0cc,
12'h0ff,
12'h0f1,
12'h0be,
12'h086,
12'h076,
12'h0b4,
12'h121,
12'h175,
12'h180,
12'h142,
12'h0ec,
12'h0c1,
12'h0e5,
12'h139,
12'h173,
12'h168,
12'h12e,
12'h0da,
12'h083,
12'h04d,
12'h058,
12'h0aa,
12'h10b,
12'h11e,
12'h0e0,
12'h0a3,
12'h08d,
12'h08e,
12'h08a,
12'h07f,
12'h05f,
12'h021,
12'hfe6,
12'hfca,
12'hfdb,
12'h000,
12'h01e,
12'h014,
12'hfd7,
12'hf80,
12'hf2a,
12'heea,
12'hec5,
12'heae,
12'he9d,
12'he92,
12'he85,
12'he73,
12'he6d,
12'he7e,
12'he91,
12'he8c,
12'he93,
12'heaa,
12'hebd,
12'hec9,
12'hebc,
12'he94,
12'he6b,
12'he5b,
12'he6c,
12'he8e,
12'hec0,
12'hf05,
12'hf4a,
12'hf61,
12'hf3c,
12'hf00,
12'hec8,
12'hea0,
12'he85,
12'he63,
12'he3f,
12'he3d,
12'he69,
12'hed6,
12'hf6f,
12'hfea,
12'h028,
12'h02d,
12'hff6,
12'hf95,
12'hf2e,
12'hedf,
12'heb0,
12'hea0,
12'heb1,
12'hee5,
12'hf35,
12'hf9b,
12'h00a,
12'h06f,
12'h0b9,
12'h0e5,
12'h0f5,
12'h0d7,
12'h07a,
12'hffd,
12'hf95,
12'hf66,
12'hf78,
12'hfbc,
12'h036,
12'h0d8,
12'h169,
12'h1c4,
12'h1ec,
12'h21c,
12'h27e,
12'h2cb,
12'h2bd,
12'h246,
12'h1a7,
12'h140,
12'h132,
12'h176,
12'h1fe,
12'h2ab,
12'h319,
12'h300,
12'h28d,
12'h22e,
12'h21d,
12'h242,
12'h27a,
12'h294,
12'h25e,
12'h1dc,
12'h163,
12'h144,
12'h170,
12'h199,
12'h18e,
12'h168,
12'h13a,
12'h10e,
12'h0e1,
12'h0d7,
12'h108,
12'h11e,
12'h0e4,
12'h07e,
12'h029,
12'h003,
12'h002,
12'h019,
12'h023,
12'hff2,
12'hf70,
12'heb8,
12'he1c,
12'hdee,
12'he3c,
12'hecc,
12'hf4e,
12'hf9a,
12'hfa2,
12'hf66,
12'hf1c,
12'hefe,
12'hf0a,
12'hf16,
12'heec,
12'he8c,
12'he29,
12'he05,
12'he27,
12'he64,
12'hea7,
12'hed2,
12'hed1,
12'head,
12'he79,
12'he4d,
12'he49,
12'he94,
12'hf16,
12'hf8c,
12'hfb5,
12'hf82,
12'hf28,
12'hedb,
12'hec2,
12'heda,
12'hf04,
12'hf45,
12'hf8a,
12'hfad,
12'hfad,
12'hfbf,
12'h000,
12'h039,
12'h044,
12'h024,
12'hfdd,
12'hf90,
12'hf75,
12'hfab,
12'h012,
12'h06f,
12'h09e,
12'h0a9,
12'h0a3,
12'h09d,
12'h09b,
12'h0c0,
12'h129,
12'h196,
12'h1c0,
12'h19c,
12'h15a,
12'h123,
12'h0fb,
12'h0f1,
12'h107,
12'h11d,
12'h11d,
12'h105,
12'h0f3,
12'h0fb,
12'h10f,
12'h11c,
12'h115,
12'h103,
12'h0e9,
12'h0cc,
12'h0ae,
12'h09e,
12'h09b,
12'h08a,
12'h079,
12'h071,
12'h069,
12'h062,
12'h053,
12'h03a,
12'h00f,
12'hfd5,
12'hfac,
12'hfaa,
12'hfbe,
12'hfc0,
12'hfb6,
12'hfa6,
12'hf82,
12'hf49,
12'hef6,
12'he93,
12'he43,
12'he15,
12'he13,
12'he39,
12'he70,
12'hea2,
12'hebe,
12'hecd,
12'hedd,
12'hede,
12'hebc,
12'he79,
12'he3a,
12'he2b,
12'he35,
12'he41,
12'he76,
12'hef0,
12'hf83,
12'hfc8,
12'hfa4,
12'hf63,
12'hf2e,
12'hef2,
12'he9a,
12'he4e,
12'he4f,
12'he9e,
12'hef0,
12'hf0f,
12'hf26,
12'hf67,
12'hfc4,
12'hfef,
12'hfbb,
12'hf5e,
12'hef9,
12'he9f,
12'he7f,
12'hebb,
12'hf45,
12'hfcf,
12'h004,
12'hff1,
12'hff6,
12'h04b,
12'h0ab,
12'h0c2,
12'h08e,
12'h031,
12'hfcc,
12'hf7a,
12'hf63,
12'hf91,
12'hfeb,
12'h041,
12'h081,
12'h0ca,
12'h12c,
12'h19e,
12'h203,
12'h24a,
12'h258,
12'h20f,
12'h180,
12'h0f7,
12'h0cf,
12'h118,
12'h1a4,
12'h22e,
12'h2a1,
12'h30d,
12'h35d,
12'h374,
12'h362,
12'h34d,
12'h311,
12'h299,
12'h212,
12'h19d,
12'h158,
12'h147,
12'h170,
12'h1c8,
12'h203,
12'h1f6,
12'h1b7,
12'h180,
12'h15f,
12'h143,
12'h12f,
12'h12f,
12'h11e,
12'h0e0,
12'h085,
12'h03a,
12'h018,
12'h00f,
12'h00f,
12'hff4,
12'hfa1,
12'hf37,
12'hef5,
12'hf04,
12'hf4e,
12'hfa1,
12'hfc8,
12'hfac,
12'hf49,
12'heb9,
12'he51,
12'he49,
12'he8d,
12'hee5,
12'hf13,
12'heff,
12'hebd,
12'he76,
12'he5c,
12'he89,
12'hece,
12'heed,
12'hed1,
12'he94,
12'he63,
12'he5b,
12'he74,
12'hea8,
12'heef,
12'hf26,
12'hf27,
12'hee7,
12'hea5,
12'heaa,
12'hee8,
12'hf2f,
12'hf57,
12'hf58,
12'hf48,
12'hf42,
12'hf5b,
12'hf9e,
12'hff9,
12'h039,
12'h012,
12'hf9a,
12'hf37,
12'hf16,
12'hf4a,
12'hfb5,
12'h01b,
12'h05a,
12'h053,
12'h01d,
12'hff5,
12'h022,
12'h097,
12'h0ff,
12'h126,
12'h112,
12'h0dd,
12'h098,
12'h071,
12'h0a0,
12'h120,
12'h196,
12'h1bb,
12'h194,
12'h14a,
12'h112,
12'h104,
12'h121,
12'h14c,
12'h160,
12'h142,
12'h0fa,
12'h0a1,
12'h056,
12'h044,
12'h07b,
12'h0d9,
12'h11e,
12'h10f,
12'h0d1,
12'h0a4,
12'h0a0,
12'h0a2,
12'h08c,
12'h078,
12'h066,
12'h046,
12'h01a,
12'hff7,
12'hffd,
12'h019,
12'h02f,
12'h023,
12'hfd9,
12'hf62,
12'hedf,
12'he75,
12'he4e,
12'he67,
12'he97,
12'heb8,
12'hec7,
12'hec9,
12'heaf,
12'he87,
12'he76,
12'he88,
12'he95,
12'he7e,
12'he63,
12'he5d,
12'he64,
12'he71,
12'he7c,
12'he90,
12'hec0,
12'heed,
12'hef4,
12'hf00,
12'hf32,
12'hf59,
12'hf32,
12'hede,
12'heab,
12'hea8,
12'heb5,
12'heb3,
12'hea5,
12'hea2,
12'hea4,
12'hec0,
12'hf14,
12'hf95,
12'h00b,
12'h01f,
12'hfbf,
12'hf26,
12'hea7,
12'he81,
12'hec2,
12'hf2e,
12'hf6f,
12'hf7e,
12'hf85,
12'hfb8,
12'h020,
12'h09e,
12'h102,
12'h123,
12'h0e5,
12'h037,
12'hf7b,
12'hf1f,
12'hf35,
12'hf96,
12'h009,
12'h075,
12'h0c2,
12'h0f0,
12'h124,
12'h180,
12'h212,
12'h2a3,
12'h2df,
12'h295,
12'h1ea,
12'h13c,
12'h0e7,
12'h122,
12'h1c9,
12'h27b,
12'h2e4,
12'h2f8,
12'h2db,
12'h2bb,
12'h2ae,
12'h2b6,
12'h2ce,
12'h2c1,
12'h26a,
12'h1dc,
12'h168,
12'h15a,
12'h19e,
12'h1e1,
12'h1f0,
12'h1c3,
12'h174,
12'h120,
12'h0f1,
12'h0f9,
12'h11b,
12'h138,
12'h11e,
12'h0b0,
12'h01b,
12'hfbf,
12'hfd3,
12'h033,
12'h090,
12'h0af,
12'h086,
12'h00c,
12'hf68,
12'hecf,
12'he69,
12'he5e,
12'he9c,
12'hef5,
12'hf33,
12'hf2d,
12'hefe,
12'hee7,
12'hf0a,
12'hf4e,
12'hf71,
12'hf48,
12'hedc,
12'he5b,
12'he04,
12'hdf8,
12'he28,
12'he85,
12'heea,
12'hf10,
12'hed8,
12'he74,
12'he3b,
12'he54,
12'heb9,
12'hf35,
12'hf8c,
12'hfac,
12'hf82,
12'hf20,
12'heae,
12'he79,
12'heb3,
12'hf20,
12'hf78,
12'hf9f,
12'hf96,
12'hf84,
12'hf9e,
12'hffc,
12'h060,
12'h073,
12'h02b,
12'hfb2,
12'hf3a,
12'hefc,
12'hf25,
12'hfaa,
12'h053,
12'h0cc,
12'h0d2,
12'h07e,
12'h022,
12'h015,
12'h067,
12'h0e8,
12'h15e,
12'h197,
12'h187,
12'h145,
12'h101,
12'h0f6,
12'h113,
12'h120,
12'h105,
12'h0c6,
12'h08c,
12'h068,
12'h069,
12'h09a,
12'h0d8,
12'h0f2,
12'h0d4,
12'h097,
12'h072,
12'h07e,
12'h09d,
12'h0ae,
12'h0ac,
12'h094,
12'h068,
12'h03c,
12'h020,
12'h019,
12'h025,
12'h018,
12'hfca,
12'hf5a,
12'hf12,
12'hf20,
12'hf78,
12'hfdf,
12'h01b,
12'h002,
12'hf8f,
12'hef4,
12'he76,
12'he43,
12'he3b,
12'he3a,
12'he2e,
12'he13,
12'he14,
12'he34,
12'he75,
12'hecd,
12'hf14,
12'hf18,
12'hece,
12'he64,
12'he28,
12'he46,
12'he7b,
12'he9b,
12'hec4,
12'hf05,
12'hf40,
12'hf43,
12'hf10,
12'hef4,
12'hf0c,
12'hf22,
12'hf04,
12'hec8,
12'hea2,
12'hea1,
12'heaf,
12'hed9,
12'hf39,
12'hfb2,
12'h006,
12'h001,
12'hfb4,
12'hf5e,
12'hf43,
12'hf64,
12'hf8c,
12'hf98,
12'hf7c,
12'hf5c,
12'hf51,
12'hf70,
12'hfdd,
12'h086,
12'h110,
12'h118,
12'h09f,
12'h00a,
12'hfba,
12'hfc0,
12'hffe,
12'h046,
12'h079,
12'h07f,
12'h078,
12'h0b7,
12'h15a,
12'h217,
12'h28e,
12'h294,
12'h22b,
12'h195,
12'h123,
12'h108,
12'h14e,
12'h1d7,
12'h25d,
12'h293,
12'h28c,
12'h29f,
12'h2e9,
12'h336,
12'h33b,
12'h2fd,
12'h2a7,
12'h242,
12'h1f4,
12'h1da,
12'h1ff,
12'h23d,
12'h250,
12'h221,
12'h1c0,
12'h151,
12'h10f,
12'h112,
12'h13b,
12'h163,
12'h15c,
12'h11d,
12'h0c8,
12'h090,
12'h097,
12'h0b5,
12'h0bb,
12'h093,
12'h041,
12'hfdd,
12'hf71,
12'hf21,
12'hf11,
12'hf2e,
12'hf4f,
12'hf4b,
12'hf2d,
12'hf0b,
12'hee9,
12'hecf,
12'hecf,
12'hef9,
12'hf29,
12'hf3d,
12'hf20,
12'heeb,
12'heb3,
12'he76,
12'he43,
12'he3c,
12'he65,
12'he8d,
12'he9b,
12'he95,
12'he89,
12'he93,
12'heb5,
12'hed5,
12'hef6,
12'hf0a,
12'hf00,
12'hee2,
12'hec2,
12'hecd,
12'hef8,
12'hf39,
12'hf71,
12'hf66,
12'hf23,
12'hee3,
12'heea,
12'hf44,
12'hfce,
12'h048,
12'h065,
12'h00c,
12'hf7e,
12'hf16,
12'hf15,
12'hf65,
12'hfd6,
12'h036,
12'h058,
12'h023,
12'hfc2,
12'hfa0,
12'h000,
12'h0b2,
12'h13a,
12'h15b,
12'h125,
12'h0c8,
12'h08c,
12'h0a2,
12'h10b,
12'h188,
12'h1b8,
12'h16d,
12'h0d7,
12'h058,
12'h04e,
12'h0b7,
12'h137,
12'h184,
12'h178,
12'h119,
12'h09b,
12'h04a,
12'h064,
12'h0cd,
12'h130,
12'h145,
12'h0fd,
12'h080,
12'h01b,
12'h010,
12'h041,
12'h083,
12'h0a1,
12'h077,
12'h026,
12'hfdc,
12'hfc5,
12'hfef,
12'h02d,
12'h04e,
12'h037,
12'hfe5,
12'hf75,
12'hf0e,
12'hecf,
12'hec7,
12'hece,
12'hebc,
12'he8e,
12'he5c,
12'he4b,
12'he6c,
12'heb4,
12'hf07,
12'hf3d,
12'hf2f,
12'hee1,
12'he8b,
12'he56,
12'he4b,
12'he62,
12'he82,
12'hea5,
12'hec4,
12'hed9,
12'hef5,
12'hf2e,
12'hf72,
12'hf81,
12'hf3a,
12'hed4,
12'he9a,
12'he88,
12'he8b,
12'he95,
12'he98,
12'he98,
12'heb3,
12'hf04,
12'hf7b,
12'hfea,
12'h018,
12'hff9,
12'hf99,
12'hf25,
12'hed8,
12'hec6,
12'hed9,
12'hee2,
12'hedc,
12'hef6,
12'hf4f,
12'hfd5,
12'h06c,
12'h0f8,
12'h141,
12'h123,
12'h0b5,
12'h02c,
12'hfc7,
12'hf96,
12'hf7e,
12'hf7a,
12'hf8c,
12'hfc7,
12'h040,
12'h0f7,
12'h1b6,
12'h22f,
12'h255,
12'h250,
12'h240,
12'h21c,
12'h1d1,
12'h167,
12'h106,
12'h0f1,
12'h13d,
12'h1c1,
12'h25c,
12'h2e8,
12'h31e,
12'h2ef,
12'h286,
12'h223,
12'h202,
12'h223,
12'h25f,
12'h274,
12'h23d,
12'h1d0,
12'h173,
12'h15e,
12'h17d,
12'h192,
12'h17a,
12'h135,
12'h0e6,
12'h0ad,
12'h0a2,
12'h0cc,
12'h103,
12'h10c,
12'h0cb,
12'h060,
12'h00a,
12'hff4,
12'h01d,
12'h058,
12'h065,
12'h020,
12'hf80,
12'hea2,
12'hdf9,
12'hdf2,
12'he78,
12'hf21,
12'hf8a,
12'hf8b,
12'hf4a,
12'hf13,
12'hf15,
12'hf49,
12'hf7d,
12'hf6f,
12'hef9,
12'he4d,
12'hdc4,
12'hd9a,
12'hdd0,
12'he3d,
12'heae,
12'hef5,
12'hf00,
12'hee1,
12'heb7,
12'heb8,
12'hef4,
12'hf44,
12'hf71,
12'hf6f,
12'hf50,
12'hf10,
12'hed6,
12'hed8,
12'hf12,
12'hf4f,
12'hf5f,
12'hf54,
12'hf67,
12'hf99,
12'hfce,
12'h003,
12'h02b,
12'h03a,
12'h026,
12'hff1,
12'hfaf,
12'hf84,
12'hf90,
12'hfd8,
12'h03e,
12'h08c,
12'h0be,
12'h0d6,
12'h0d9,
12'h0d1,
12'h0ba,
12'h0b6,
12'h0e9,
12'h133,
12'h164,
12'h164,
12'h139,
12'h101,
12'h0d6,
12'h0d3,
12'h0fc,
12'h134,
12'h14f,
12'h129,
12'h0c7,
12'h078,
12'h06f,
12'h08c,
12'h0c1,
12'h10f,
12'h130,
12'h102,
12'h0be,
12'h08e,
12'h088,
12'h090,
12'h08f,
12'h074,
12'h039,
12'hffe,
12'hfcc,
12'hfb0,
12'hfb3,
12'hfd6,
12'hff7,
12'h001,
12'hff9,
12'hfd5,
12'hfbb,
12'hfa9,
12'hf87,
12'hf3e,
12'hed4,
12'he73,
12'he1f,
12'hdea,
12'hdef,
12'he30,
12'he90,
12'hedc,
12'hef9,
12'hf00,
12'hf04,
12'heed,
12'heb1,
12'he7c,
12'he6c,
12'he6b,
12'he51,
12'he33,
12'he6a,
12'hefb,
12'hf90,
12'hfd7,
12'hfbb,
12'hf87,
12'hf58,
12'hf0c,
12'heb3,
12'he81,
12'he96,
12'hecc,
12'heeb,
12'heec,
12'heea,
12'hf1c,
12'hf73,
12'hfb1,
12'hfb9,
12'hf82,
12'hf2c,
12'hed6,
12'heaf,
12'hed7,
12'hf45,
12'hfd0,
12'h026,
12'h034,
12'h03f,
12'h063,
12'h07e,
12'h07e,
12'h05c,
12'h01d,
12'hfc7,
12'hf79,
12'hf70,
12'hfc8,
12'h04e,
12'h0b8,
12'h107,
12'h153,
12'h186,
12'h189,
12'h186,
12'h19b,
12'h1af,
12'h190,
12'h13b,
12'h0ec,
12'h0ec,
12'h150,
12'h1e2,
12'h270,
12'h2e5,
12'h335,
12'h339,
12'h2ff,
12'h2d7,
12'h2d2,
12'h2bc,
12'h26f,
12'h204,
12'h197,
12'h148,
12'h13c,
12'h17b,
12'h1e6,
12'h239,
12'h228,
12'h1c5,
12'h172,
12'h159,
12'h16c,
12'h180,
12'h16a,
12'h116,
12'h09a,
12'h03c,
12'h01c,
12'h033,
12'h06a,
12'h084,
12'h049,
12'hfba,
12'hf2f,
12'hef0,
12'hf11,
12'hf78,
12'hfcf,
12'hfcc,
12'hf5a,
12'hec1,
12'he5f,
12'he64,
12'hebe,
12'hf0f,
12'hf23,
12'heff,
12'hebf,
12'he88,
12'he7d,
12'heac,
12'hef0,
12'hf13,
12'heee,
12'he7e,
12'he1e,
12'he20,
12'he74,
12'hed5,
12'hf0b,
12'hf0e,
12'hef0,
12'hecb,
12'heb4,
12'hec0,
12'hef4,
12'hf2c,
12'hf41,
12'hf22,
12'hefa,
12'hf02,
12'hf36,
12'hf8e,
12'hfd8,
12'hffd,
12'hfec,
12'hf95,
12'hf3f,
12'hf1f,
12'hf48,
12'hf9d,
12'hfe1,
12'h00b,
12'h01c,
12'h00e,
12'hffa,
12'h009,
12'h04a,
12'h08e,
12'h0ac,
12'h09a,
12'h089,
12'h0a8,
12'h0cd,
12'h0db,
12'h0f0,
12'h11f,
12'h147,
12'h149,
12'h135,
12'h122,
12'h114,
12'h104,
12'h0f9,
12'h0fa,
12'h109,
12'h109,
12'h0e2,
12'h0ab,
12'h067,
12'h033,
12'h03d,
12'h088,
12'h0d6,
12'h0f0,
12'h0d5,
12'h0a8,
12'h08e,
12'h07c,
12'h072,
12'h06e,
12'h064,
12'h042,
12'hff9,
12'hfb7,
12'hfa7,
12'hfbf,
12'hfe2,
12'hfe8,
12'hfc6,
12'hf76,
12'hef4,
12'he7d,
12'he49,
12'he60,
12'he95,
12'heae,
12'hea6,
12'he9a,
12'he96,
12'he9d,
12'hebd,
12'hee9,
12'hefb,
12'hed5,
12'he97,
12'he68,
12'he5a,
12'he6d,
12'he94,
12'hebb,
12'hedc,
12'hee2,
12'hedb,
12'hef7,
12'hf3a,
12'hf81,
12'hf8d,
12'hf5a,
12'hf17,
12'hee3,
12'hebd,
12'he9a,
12'hea3,
12'hec4,
12'heda,
12'hede,
12'hee4,
12'hf38,
12'hfb9,
12'h009,
12'hfe9,
12'hf6c,
12'hedc,
12'he79,
12'he76,
12'hec3,
12'hf3e,
12'hfbc,
12'h004,
12'h024,
12'h047,
12'h08f,
12'h0e4,
12'h105,
12'h0d5,
12'h044,
12'hf93,
12'hf1a,
12'hf0c,
12'hf69,
12'hff1,
12'h088,
12'h11f,
12'h196,
12'h1c7,
12'h1bc,
12'h1d1,
12'h229,
12'h27c,
12'h265,
12'h1d6,
12'h133,
12'h0ec,
12'h125,
12'h1bf,
12'h276,
12'h306,
12'h329,
12'h2d6,
12'h257,
12'h21f,
12'h23f,
12'h282,
12'h2b3,
12'h293,
12'h215,
12'h16f,
12'h119,
12'h14d,
12'h1d1,
12'h22c,
12'h21b,
12'h1be,
12'h14a,
12'h0e3,
12'h0a1,
12'h0a5,
12'h0ed,
12'h120,
12'h0e9,
12'h069,
12'hffb,
12'hfe9,
12'h024,
12'h081,
12'h0be,
12'h08e,
12'hff2,
12'hf24,
12'he86,
12'he42,
12'he61,
12'hecd,
12'hf4a,
12'hfa2,
12'hfa2,
12'hf5e,
12'hf1e,
12'hf19,
12'hf48,
12'hf64,
12'hf2e,
12'hea9,
12'he20,
12'hdcd,
12'hdc7,
12'he1b,
12'heae,
12'hf4b,
12'hf99,
12'hf6a,
12'hefa,
12'he9b,
12'he85,
12'heb9,
12'hf13,
12'hf63,
12'hf77,
12'hf47,
12'heef,
12'hea9,
12'hea6,
12'heea,
12'hf53,
12'hfac,
12'hfde,
12'hfdf,
12'hfbb,
12'hfbc,
12'h008,
12'h06a,
12'h08d,
12'h053,
12'hfd9,
12'hf58,
12'hf17,
12'hf3a,
12'hfb7,
12'h062,
12'h0eb,
12'h111,
12'h0e0,
12'h08e,
12'h064,
12'h096,
12'h109,
12'h16e,
12'h183,
12'h154,
12'h115,
12'h0ef,
12'h0ee,
12'h112,
12'h148,
12'h164,
12'h148,
12'h0fe,
12'h0a2,
12'h05a,
12'h044,
12'h068,
12'h0b3,
12'h0f7,
12'h104,
12'h0d8,
12'h0b6,
12'h0b2,
12'h0a4,
12'h081,
12'h056,
12'h047,
12'h036,
12'h00c,
12'hfe6,
12'hfdf,
12'hff2,
12'hff0,
12'hfcb,
12'hfa5,
12'hf98,
12'hfa3,
12'hfaa,
12'hfb7,
12'hfb1,
12'hf76,
12'hf0b,
12'he8a,
12'he3a,
12'he23,
12'he2f,
12'he45,
12'he54,
12'he66,
12'he81,
12'heae,
12'hee3,
12'hf10,
12'hf12,
12'hed4,
12'he85,
12'he5d,
12'he5c,
12'he59,
12'he5d,
12'he9e,
12'hf0a,
12'hf5c,
12'hf6d,
12'hf59,
12'hf4f,
12'hf3a,
12'hf00,
12'hebb,
12'he91,
12'he87,
12'he87,
12'he80,
12'hea2,
12'hf16,
12'hf9a,
12'hfd7,
12'hfb7,
12'hf63,
12'hf17,
12'hef3,
12'hf06,
12'hf3d,
12'hf74,
12'hf91,
12'hf92,
12'hf9b,
12'hfc0,
12'hff5,
12'h02e,
12'h058,
12'h04e,
12'hfff,
12'hf8e,
12'hf53,
12'hf78,
12'hfdb,
12'h048,
12'h08b,
12'h097,
12'h09c,
12'h0ce,
12'h135,
12'h1b0,
12'h207,
12'h218,
12'h1d2,
12'h15f,
12'h10c,
12'h107,
12'h15e,
12'h1e5,
12'h25c,
12'h28b,
12'h290,
12'h2ad,
12'h2e5,
12'h30c,
12'h2fd,
12'h2c1,
12'h26b,
12'h214,
12'h1c3,
12'h188,
12'h18a,
12'h1d3,
12'h21f,
12'h225,
12'h1e3,
12'h181,
12'h13b,
12'h11e,
12'h120,
12'h132,
12'h129,
12'h0f2,
12'h09f,
12'h071,
12'h084,
12'h0b2,
12'h0cb,
12'h0a4,
12'h04a,
12'hfbc,
12'hf22,
12'hede,
12'hefd,
12'hf53,
12'hf8c,
12'hf8f,
12'hf7b,
12'hf4a,
12'hf06,
12'hed2,
12'hede,
12'hf15,
12'hf38,
12'hf32,
12'hef4,
12'heb2,
12'he8d,
12'he7f,
12'hea5,
12'hee5,
12'hf07,
12'hee1,
12'he8d,
12'he5b,
12'he68,
12'heaa,
12'hee8,
12'hf12,
12'hf17,
12'hef3,
12'hec7,
12'heb0,
12'hed0,
12'hf05,
12'hf22,
12'hf2c,
12'hf33,
12'hf3a,
12'hf48,
12'hf73,
12'hfb3,
12'hff8,
12'h01a,
12'hff6,
12'hfa0,
12'hf45,
12'hf10,
12'hf13,
12'hf45,
12'hf97,
12'hfe7,
12'h01b,
12'h028,
12'h011,
12'h00a,
12'h033,
12'h089,
12'h0df,
12'h10d,
12'h117,
12'h0fa,
12'h0cd,
12'h0c3,
12'h0f3,
12'h145,
12'h178,
12'h15b,
12'h102,
12'h0ac,
12'h086,
12'h09b,
12'h0db,
12'h11f,
12'h135,
12'h106,
12'h0a7,
12'h049,
12'h039,
12'h08b,
12'h100,
12'h140,
12'h119,
12'h0b6,
12'h05a,
12'h027,
12'h019,
12'h02c,
12'h059,
12'h071,
12'h052,
12'h006,
12'hfc4,
12'hfc0,
12'hff0,
12'h022,
12'h021,
12'hfea,
12'hf89,
12'hf10,
12'heb5,
12'he9c,
12'heca,
12'hf05,
12'hf20,
12'hf10,
12'hed4,
12'he8a,
12'he64,
12'he84,
12'hed0,
12'hf0e,
12'hf0b,
12'heca,
12'he84,
12'he5f,
12'he59,
12'he91,
12'hee7,
12'hf28,
12'hf36,
12'hf1a,
12'hf16,
12'hf3b,
12'hf70,
12'hf84,
12'hf5e,
12'hf23,
12'heef,
12'hec3,
12'hea2,
12'he8c,
12'he89,
12'heb1,
12'hf14,
12'hf96,
12'hffd,
12'h03b,
12'h049,
12'h00d,
12'hf9a,
12'hf31,
12'hf01,
12'heff,
12'hf05,
12'hef2,
12'heeb,
12'hf29,
12'hf9f,
12'h038,
12'h0d3,
12'h137,
12'h13b,
12'h0e3,
12'h055,
12'hfce,
12'hf89,
12'hf9a,
12'hfd4,
12'hffe,
12'h015,
12'h03e,
12'h09b,
12'h138,
12'h1ee,
12'h274,
12'h2af,
12'h2ad,
12'h273,
12'h207,
12'h193,
12'h148,
12'h13f,
12'h174,
12'h1b9,
12'h1fc,
12'h254,
12'h2a5,
12'h2bd,
12'h29b,
12'h265,
12'h243,
12'h240,
12'h24b,
12'h243,
12'h211,
12'h1c4,
12'h185,
12'h16d,
12'h174,
12'h171,
12'h14e,
12'h11b,
12'h101,
12'h0ea,
12'h0b9,
12'h095,
12'h08b,
12'h082,
12'h072,
12'h05c,
12'h048,
12'h048,
12'h04c,
12'h041,
12'h020,
12'hfe3,
12'hf87,
12'hf08,
12'he70,
12'he12,
12'he28,
12'he92,
12'hf1a,
12'hf7c,
12'hfa3,
12'hf99,
12'hf76,
12'hf5d,
12'hf50,
12'hf42,
12'hf13,
12'hebd,
12'he60,
12'he17,
12'he0b,
12'he46,
12'he9d,
12'hee8,
12'hf0b,
12'hf00,
12'hed0,
12'he9c,
12'he89,
12'heaf,
12'hf08,
12'hf68,
12'hf92,
12'hf6b,
12'hf02,
12'heae,
12'heb9,
12'hf03,
12'hf54,
12'hf83,
12'hf9a,
12'hfa5,
12'hfac,
12'hfc2,
12'hfed,
12'h003,
12'hfee,
12'hfb9,
12'hf79,
12'hf4f,
12'hf64,
12'hfc2,
12'h03b,
12'h092,
12'h09a,
12'h074,
12'h059,
12'h066,
12'h088,
12'h0bf,
12'h115,
12'h166,
12'h18f,
12'h174,
12'h139,
12'h114,
12'h0fe,
12'h0ee,
12'h0e8,
12'h0fb,
12'h118,
12'h113,
12'h0f6,
12'h0db,
12'h0c3,
12'h0ae,
12'h0a4,
12'h0ae,
12'h0c1,
12'h0d4,
12'h0e1,
12'h0d5,
12'h0b4,
12'h07f,
12'h049,
12'h03a,
12'h042,
12'h043,
12'h029,
12'hff1,
12'hfab,
12'hf7b,
12'hf83,
12'hfbb,
12'hff6,
12'h016,
12'h009,
12'hfc7,
12'hf65,
12'hf12,
12'heeb,
12'hecf,
12'hea3,
12'he59,
12'he1e,
12'he21,
12'he59,
12'hea0,
12'hecb,
12'hed8,
12'hed5,
12'hec5,
12'he9f,
12'he6f,
12'he61,
12'he7b,
12'he9f,
12'hea5,
12'he97,
12'hebd,
12'hf16,
12'hf68,
12'hf87,
12'hf80,
12'hf6c,
12'hf31,
12'hed9,
12'he89,
12'he6c,
12'he91,
12'hecd,
12'heef,
12'heec,
12'hefe,
12'hf41,
12'hf83,
12'hf9a,
12'hf7c,
12'hf3a,
12'hed9,
12'he91,
12'hea2,
12'hf11,
12'hf9d,
12'hfe5,
12'hfea,
12'hff8,
12'h03f,
12'h096,
12'h0b1,
12'h082,
12'h024,
12'hfba,
12'hf5b,
12'hf40,
12'hf88,
12'h00a,
12'h079,
12'h0b8,
12'h0f2,
12'h130,
12'h16d,
12'h19b,
12'h1b0,
12'h1a9,
12'h176,
12'h121,
12'h0d3,
12'h0dd,
12'h168,
12'h219,
12'h295,
12'h2e1,
12'h319,
12'h338,
12'h32a,
12'h308,
12'h2f8,
12'h2e4,
12'h2a9,
12'h250,
12'h1fc,
12'h1b3,
12'h187,
12'h195,
12'h1d5,
12'h20b,
12'h1f8,
12'h1ae,
12'h174,
12'h164,
12'h167,
12'h16c,
12'h15b,
12'h12c,
12'h0dc,
12'h083,
12'h052,
12'h053,
12'h076,
12'h08e,
12'h06d,
12'h00f,
12'hf98,
12'hf39,
12'hf20,
12'hf50,
12'hf98,
12'hfbe,
12'hf98,
12'hf30,
12'hec2,
12'he98,
12'hece,
12'hf21,
12'hf56,
12'hf62,
12'hf2e,
12'hed8,
12'he88,
12'he68,
12'he98,
12'hedf,
12'hf04,
12'hee0,
12'he8e,
12'he59,
12'he5a,
12'he80,
12'heb7,
12'heec,
12'hf0f,
12'hf1b,
12'hf0a,
12'hee7,
12'hed3,
12'hee0,
12'hefa,
12'hf03,
12'hef1,
12'hede,
12'heee,
12'hf2c,
12'hf7e,
12'hfd1,
12'h014,
12'h014,
12'hfb9,
12'hf41,
12'hf00,
12'hf14,
12'hf52,
12'hfa0,
12'hfe2,
12'hff4,
12'hfe0,
12'hfd7,
12'h003,
12'h061,
12'h0bb,
12'h0de,
12'h0c6,
12'h09a,
12'h076,
12'h06f,
12'h09b,
12'h0fb,
12'h166,
12'h186,
12'h146,
12'h0eb,
12'h0ad,
12'h0b8,
12'h100,
12'h145,
12'h168,
12'h152,
12'h103,
12'h093,
12'h03b,
12'h02e,
12'h069,
12'h0c8,
12'h100,
12'h0f9,
12'h0c0,
12'h089,
12'h08b,
12'h0a5,
12'h0b2,
12'h09d,
12'h05b,
12'h007,
12'hfc6,
12'hfb2,
12'hfd0,
12'h00b,
12'h036,
12'h041,
12'h01b,
12'hfb9,
12'hf32,
12'heae,
12'he6d,
12'he6f,
12'he86,
12'he9f,
12'hea4,
12'hea3,
12'hea7,
12'heac,
12'hec2,
12'heda,
12'hef0,
12'heee,
12'heca,
12'heb9,
12'heb4,
12'head,
12'heab,
12'hebc,
12'hede,
12'heed,
12'hee8,
12'heec,
12'hf06,
12'hf18,
12'hf05,
12'hedd,
12'hecd,
12'heda,
12'hed4,
12'he9a,
12'he4c,
12'he2b,
12'he58,
12'heba,
12'hf27,
12'hf92,
12'hfe5,
12'h000,
12'hfda,
12'hf95,
12'hf60,
12'hf2a,
12'hef1,
12'hec4,
12'hebc,
12'hee4,
12'hf2f,
12'hf8c,
12'hfec,
12'h054,
12'h0b2,
12'h0ec,
12'h0ed,
12'h09f,
12'h015,
12'hf84,
12'hf29,
12'hf2d,
12'hf79,
12'hfdd,
12'h064,
12'h10d,
12'h1a2,
12'h1f8,
12'h20d,
12'h22c,
12'h26e,
12'h29a,
12'h26b,
12'h1e1,
12'h164,
12'h144,
12'h187,
12'h1f4,
12'h274,
12'h2e4,
12'h2e9,
12'h29b,
12'h242,
12'h21c,
12'h245,
12'h290,
12'h2d8,
12'h2d9,
12'h27b,
12'h203,
12'h19e,
12'h185,
12'h1a3,
12'h1b0,
12'h198,
12'h159,
12'h12e,
12'h124,
12'h12f,
12'h156,
12'h16c,
12'h148,
12'h0e3,
12'h06e,
12'h02d,
12'h039,
12'h079,
12'h0ac,
12'h096,
12'h022,
12'hf60,
12'he88,
12'hdf5,
12'hdee,
12'he54,
12'hed4,
12'hf4f,
12'hfa7,
12'hfc6,
12'hfaa,
12'hf80,
12'hf72,
12'hf5a,
12'hf16,
12'he9b,
12'he15,
12'hdc8,
12'hdd6,
12'he31,
12'he95,
12'heee,
12'hf23,
12'hf1f,
12'hee5,
12'he85,
12'he3d,
12'he31,
12'he6f,
12'heea,
12'hf68,
12'hfb0,
12'hfa1,
12'hf42,
12'hee0,
12'heba,
12'heca,
12'hefe,
12'hf3e,
12'hf73,
12'hf8a,
12'hf8d,
12'hfac,
12'hfee,
12'h022,
12'h018,
12'hfc9,
12'hf5d,
12'hf18,
12'hf29,
12'hf8a,
12'h001,
12'h065,
12'h0a3,
12'h0b7,
12'h095,
12'h057,
12'h02e,
12'h046,
12'h0c4,
12'h153,
12'h19d,
12'h188,
12'h139,
12'h0f6,
12'h0cb,
12'h0c6,
12'h0dc,
12'h0ed,
12'h0ea,
12'h0c7,
12'h0a7,
12'h0a4,
12'h0cc,
12'h111,
12'h145,
12'h140,
12'h0fa,
12'h0ab,
12'h08a,
12'h098,
12'h0ab,
12'h096,
12'h079,
12'h066,
12'h04b,
12'h034,
12'h02e,
12'h033,
12'h020,
12'hfe5,
12'hf9d,
12'hf6d,
12'hf71,
12'hf97,
12'hfbe,
12'hfcb,
12'hfae,
12'hf6f,
12'hf1c,
12'hecf,
12'he99,
12'he72,
12'he65,
12'he71,
12'he89,
12'hea8,
12'hec5,
12'hee4,
12'hf04,
12'hef8,
12'heb0,
12'he47,
12'he0d,
12'he32,
12'he75,
12'hea9,
12'hede,
12'hf32,
12'hf83,
12'hf84,
12'hf45,
12'hf07,
12'hefa,
12'hef5,
12'heb5,
12'he6a,
12'he65,
12'hea0,
12'hee9,
12'hf21,
12'hf6c,
12'hfdb,
12'h01f,
12'hff0,
12'hf77,
12'hf23,
12'hef3,
12'hedd,
12'heeb,
12'hf13,
12'hf40,
12'hf50,
12'hf51,
12'hf70,
12'hfcc,
12'h041,
12'h08d,
12'h093,
12'h04e,
12'hfdb,
12'hf70,
12'hf52,
12'hfa2,
12'h020,
12'h07f,
12'h094,
12'h083,
12'h0ab,
12'h119,
12'h1a9,
12'h21e,
12'h24c,
12'h230,
12'h1b0,
12'h10b,
12'h09f,
12'h0b3,
12'h14c,
12'h201,
12'h27b,
12'h2a8,
12'h2c2,
12'h2f7,
12'h323,
12'h329,
12'h308,
12'h2c1,
12'h25b,
12'h1ef,
12'h1a8,
12'h1a5,
12'h1e0,
12'h226,
12'h23e,
12'h215,
12'h1bd,
12'h165,
12'h12b,
12'h122,
12'h144,
12'h15e,
12'h147,
12'h0fc,
12'h0a4,
12'h06f,
12'h06d,
12'h087,
12'h08c,
12'h059,
12'h004,
12'hf8e,
12'hf11,
12'hed8,
12'hefa,
12'hf4b,
12'hf7d,
12'hf78,
12'hf3f,
12'heca,
12'he5c,
12'he3f,
12'he7d,
12'hed3,
12'hef5,
12'heeb,
12'hec1,
12'he9a,
12'he84,
12'he77,
12'he96,
12'hebf,
12'hec5,
12'he94,
12'he51,
12'he3b,
12'he4b,
12'he78,
12'hea7,
12'hecf,
12'hef4,
12'hf01,
12'hee7,
12'hec4,
12'heba,
12'hec4,
12'hee6,
12'hf18,
12'hf3d,
12'hf45,
12'hf43,
12'hf59,
12'hf9e,
12'h001,
12'h04d,
12'h044,
12'hfe1,
12'hf68,
12'hf28,
12'hf37,
12'hf7d,
12'hfda,
12'h026,
12'h039,
12'h01f,
12'h013,
12'h043,
12'h0b4,
12'h12f,
12'h16e,
12'h160,
12'h118,
12'h0cc,
12'h0a8,
12'h0c5,
12'h124,
12'h185,
12'h1ab,
12'h17b,
12'h113,
12'h0b5,
12'h0a7,
12'h0fc,
12'h15c,
12'h18e,
12'h189,
12'h14c,
12'h0ee,
12'h092,
12'h081,
12'h0c7,
12'h125,
12'h152,
12'h125,
12'h0c7,
12'h070,
12'h04f,
12'h063,
12'h095,
12'h0cc,
12'h0c8,
12'h079,
12'h020,
12'hfeb,
12'hfe3,
12'h000,
12'h020,
12'h023,
12'hfe6,
12'hf72,
12'hef3,
12'hea7,
12'heb7,
12'hee1,
12'heed,
12'hed5,
12'hea9,
12'he83,
12'he71,
12'he88,
12'heb7,
12'hed9,
12'heda,
12'heb3,
12'he74,
12'he51,
12'he45,
12'he3f,
12'he55,
12'he82,
12'heae,
12'hebf,
12'heba,
12'hec3,
12'heef,
12'hf0c,
12'heec,
12'hea4,
12'he7c,
12'he85,
12'he84,
12'he64,
12'he42,
12'he50,
12'he9a,
12'hefd,
12'hf53,
12'hfa0,
12'hfe4,
12'hffb,
12'hfd9,
12'hf94,
12'hf49,
12'hf03,
12'hed7,
12'heb7,
12'he9d,
12'heaf,
12'hf02,
12'hf93,
12'h03b,
12'h0c9,
12'h10d,
12'h109,
12'h0da,
12'h08a,
12'h033,
12'hff9,
12'hfe0,
12'hfda,
12'hfd7,
12'hfe9,
12'h02f,
12'h0c2,
12'h185,
12'h228,
12'h27a,
12'h298,
12'h2b0,
12'h2ba,
12'h28f,
12'h21e,
12'h1a2,
12'h16e,
12'h198,
12'h1f1,
12'h253,
12'h2bb,
12'h2fb,
12'h2fb,
12'h2bd,
12'h26b,
12'h246,
12'h250,
12'h269,
12'h25e,
12'h22a,
12'h1eb,
12'h1b7,
12'h1a3,
12'h19e,
12'h187,
12'h167,
12'h14b,
12'h130,
12'h111,
12'h0f7,
12'h0e2,
12'h0ca,
12'h0b2,
12'h090,
12'h072,
12'h05a,
12'h038,
12'h010,
12'hfe8,
12'hfbc,
12'hf72,
12'hf0d,
12'hea6,
12'he49,
12'he14,
12'he1a,
12'he6b,
12'hef0,
12'hf5a,
12'hf84,
12'hf63,
12'hf13,
12'hedf,
12'hed3,
12'hed4,
12'hec1,
12'he83,
12'he35,
12'he0c,
12'he1b,
12'he45,
12'he86,
12'hed6,
12'hefb,
12'hed3,
12'he88,
12'he57,
12'he62,
12'hea2,
12'hef8,
12'hf43,
12'hf6a,
12'hf64,
12'hf31,
12'hef1,
12'hedd,
12'hf04,
12'hf3d,
12'hf72,
12'hfa1,
12'hfad,
12'hf9c,
12'hfa2,
12'hfcc,
12'h002,
12'h02d,
12'h034,
12'h008,
12'hfd4,
12'hfd5,
12'h00e,
12'h066,
12'h0a7,
12'h0bc,
12'h0bf,
12'h0ad,
12'h09d,
12'h0b1,
12'h0fc,
12'h15e,
12'h19f,
12'h1b1,
12'h193,
12'h151,
12'h10d,
12'h0de,
12'h0d4,
12'h0ef,
12'h118,
12'h13b,
12'h144,
12'h130,
12'h10e,
12'h0fb,
12'h0f7,
12'h0ed,
12'h0ef,
12'h0f0,
12'h0e9,
12'h0d6,
12'h0ae,
12'h080,
12'h060,
12'h061,
12'h06b,
12'h068,
12'h05b,
12'h03a,
12'h009,
12'hfdb,
12'hfba,
12'hfb0,
12'hfad,
12'hfa8,
12'hf99,
12'hf85,
12'hf79,
12'hf5d,
12'hf16,
12'hebd,
12'he71,
12'he35,
12'he1f,
12'he3d,
12'he6e,
12'he96,
12'hea6,
12'he98,
12'he81,
12'he6c,
12'he4f,
12'he2a,
12'he1a,
12'he34,
12'he58,
12'he6d,
12'he76,
12'he8c,
12'hece,
12'hf09,
12'hf0b,
12'hedb,
12'hea8,
12'he92,
12'he70,
12'he34,
12'he06,
12'he0d,
12'he53,
12'he98,
12'hec5,
12'hef4,
12'hf3c,
12'hf8e,
12'hfa0,
12'hf7c,
12'hf4c,
12'hf10,
12'hed0,
12'head,
12'hecf,
12'hf1d,
12'hf63,
12'hf84,
12'hf94,
12'hfc4,
12'h028,
12'h091,
12'h0b7,
12'h094,
12'h039,
12'hfcb,
12'hf64,
12'hf39,
12'hf6b,
12'hfd1,
12'h033,
12'h08b,
12'h0f0,
12'h154,
12'h1a7,
12'h1da,
12'h1fc,
12'h20c,
12'h1da,
12'h17b,
12'h134,
12'h14c,
12'h1ce,
12'h268,
12'h2e1,
12'h325,
12'h33a,
12'h333,
12'h309,
12'h2ea,
12'h2f2,
12'h2fb,
12'h2e3,
12'h298,
12'h22a,
12'h1c2,
12'h194,
12'h1b2,
12'h1f2,
12'h20d,
12'h1d9,
12'h18f,
12'h15c,
12'h14a,
12'h165,
12'h18c,
12'h1a0,
12'h186,
12'h137,
12'h0dc,
12'h099,
12'h08c,
12'h0a3,
12'h0a8,
12'h07e,
12'h00c,
12'hf75,
12'hf16,
12'hf16,
12'hf5d,
12'hfb3,
12'hfd7,
12'hfb0,
12'hf36,
12'heab,
12'he6b,
12'hea2,
12'hf2b,
12'hf94,
12'hf93,
12'hf31,
12'heb0,
12'he4c,
12'he3a,
12'he8b,
12'hef0,
12'hf08,
12'hece,
12'he88,
12'he60,
12'he64,
12'he91,
12'hed6,
12'hf1a,
12'hf36,
12'hf1e,
12'hef4,
12'heed,
12'hf1a,
12'hf63,
12'hf8e,
12'hf7b,
12'hf4e,
12'hf29,
12'hf1b,
12'hf2a,
12'hf67,
12'hfc3,
12'h010,
12'h015,
12'hfc6,
12'hf78,
12'hf62,
12'hf89,
12'hfd2,
12'h019,
12'h03a,
12'h023,
12'hff7,
12'hff8,
12'h03b,
12'h0a2,
12'h101,
12'h123,
12'h111,
12'h0e9,
12'h0c0,
12'h0a0,
12'h09f,
12'h0c5,
12'h0ff,
12'h12c,
12'h124,
12'h0f6,
12'h0d0,
12'h0cf,
12'h0e7,
12'h0f9,
12'h0f2,
12'h0d3,
12'h0a1,
12'h062,
12'h034,
12'h049,
12'h0a6,
12'h0f9,
12'h101,
12'h0c4,
12'h073,
12'h039,
12'h01c,
12'h013,
12'h023,
12'h040,
12'h048,
12'h025,
12'hfe5,
12'hfb6,
12'hfa7,
12'hfa3,
12'hfa0,
12'hf9e,
12'hf81,
12'hf2a,
12'heab,
12'he53,
12'he48,
12'he67,
12'he89,
12'he8f,
12'he86,
12'he7a,
12'he6f,
12'he6a,
12'he7c,
12'heae,
12'hee3,
12'hedb,
12'he98,
12'he59,
12'he33,
12'he38,
12'he63,
12'heac,
12'hef8,
12'hf13,
12'heff,
12'hef6,
12'hf1c,
12'hf45,
12'hf4b,
12'hf44,
12'hf51,
12'hf53,
12'hf2a,
12'hef1,
12'hed6,
12'hf05,
12'hf59,
12'hf96,
12'hf9f,
12'hf77,
12'hf52,
12'hf42,
12'hf30,
12'hf16,
12'hefd,
12'hef0,
12'hee5,
12'hede,
12'hf0d,
12'hf8a,
12'h02c,
12'h0ba,
12'h119,
12'h149,
12'h148,
12'h10e,
12'h0ab,
12'h040,
12'hfde,
12'hf94,
12'hf79,
12'hf9c,
12'h008,
12'h097,
12'h12d,
12'h1d0,
12'h241,
12'h251,
12'h21b,
12'h1f0,
12'h1f4,
12'h1ec,
12'h19c,
12'h118,
12'h0b5,
12'h0b0,
12'h120,
12'h1e9,
12'h2c5,
12'h36a,
12'h3a7,
12'h37c,
12'h302,
12'h287,
12'h231,
12'h1f3,
12'h1c8,
12'h19d,
12'h16a,
12'h134,
12'h125,
12'h161,
12'h1c4,
12'h204,
12'h203,
12'h1d3,
12'h175,
12'h0f4,
12'h07a,
12'h028,
12'hffa,
12'hfd0,
12'hfa2,
12'hf8b,
12'hf99,
12'hfd1,
12'h02b,
12'h08d,
12'h0c2,
12'h082,
12'hfe3,
12'hf22,
12'he6b,
12'he05,
12'he0b,
12'he6e,
12'hef3,
12'hf4e,
12'hf60,
12'hf34,
12'hf07,
12'hf07,
12'hf32,
12'hf46,
12'hf09,
12'he9e,
12'he3d,
12'he0e,
12'he1c,
12'he54,
12'hea2,
12'heea,
12'hf12,
12'hf14,
12'hefc,
12'heea,
12'hefd,
12'hf32,
12'hf76,
12'hfa1,
12'hf90,
12'hf39,
12'hec2,
12'he7d,
12'he91,
12'hed9,
12'hf33,
12'hfa3,
12'h00a,
12'h030,
12'h013,
12'hffc,
12'h007,
12'h008,
12'hfe3,
12'hfa4,
12'hf63,
12'hf45,
12'hf72,
12'hfdc,
12'h060,
12'h0c9,
12'h0fb,
12'h10f,
12'h104,
12'h0db,
12'h0b1,
12'h0b3,
12'h0e7,
12'h128,
12'h148,
12'h148,
12'h13b,
12'h12a,
12'h116,
12'h10b,
12'h11d,
12'h148,
12'h161,
12'h145,
12'h101,
12'h0b4,
12'h086,
12'h064,
12'h054,
12'h075,
12'h09c,
12'h0b2,
12'h0bd,
12'h0c6,
12'h0d5,
12'h0f1,
12'h107,
12'h0fd,
12'h0c1,
12'h068,
12'h002,
12'hf92,
12'hf46,
12'hf45,
12'hf86,
12'hfd8,
12'h00a,
12'h015,
12'h003,
12'hfde,
12'hfad,
12'hf6d,
12'hf12,
12'heab,
12'he48,
12'he02,
12'hdf3,
12'he0c,
12'he41,
12'he83,
12'heac,
12'heb8,
12'heb9,
12'hebe,
12'hec5,
12'hec4,
12'hebf,
12'heab,
12'he84,
12'he5a,
12'he58,
12'he89,
12'hec9,
12'hee6,
12'hed7,
12'hed2,
12'hee9,
12'hee8,
12'hebe,
12'he9b,
12'he9e,
12'hea1,
12'he72,
12'he45,
12'he59,
12'head,
12'hefa,
12'hf0f,
12'hf12,
12'hf17,
12'hf1f,
12'hf2e,
12'hf4e,
12'hf88,
12'hfbb,
12'hfc1,
12'hfaf,
12'hfba,
12'hff8,
12'h039,
12'h047,
12'h00e,
12'hfa7,
12'hf5e,
12'hf4d,
12'hf86,
12'h007,
12'h078,
12'h0ad,
12'h0cb,
12'h0f0,
12'h11b,
12'h133,
12'h132,
12'h132,
12'h13a,
12'h11b,
12'h0c9,
12'h0a5,
12'h0f3,
12'h1a7,
12'h279,
12'h314,
12'h367,
12'h384,
12'h37a,
12'h33d,
12'h2dc,
12'h282,
12'h234,
12'h1f3,
12'h1cc,
12'h1c7,
12'h1df,
12'h1fd,
12'h21b,
12'h242,
12'h255,
12'h230,
12'h1d7,
12'h186,
12'h159,
12'h142,
12'h139,
12'h12a,
12'h113,
12'h0f0,
12'h0b8,
12'h09b,
12'h0b1,
12'h0c8,
12'h0b4,
12'h07d,
12'h03d,
12'hffd,
12'hfcf,
12'hfbc,
12'hfb5,
12'hfa8,
12'hf90,
12'hf77,
12'hf53,
12'hf33,
12'hf30,
12'hf51,
12'hf77,
12'hf6e,
12'hf31,
12'hef1,
12'heca,
12'heab,
12'he95,
12'he98,
12'hea9,
12'heb6,
12'hec3,
12'hecb,
12'hed7,
12'hedf,
12'hecb,
12'head,
12'he92,
12'he8c,
12'he94,
12'he93,
12'hea7,
12'hee7,
12'hf28,
12'hf3f,
12'hf2a,
12'hf09,
12'hf05,
12'hf25,
12'hf59,
12'hf8d,
12'hfae,
12'hfab,
12'hf90,
12'hf75,
12'hf68,
12'hf75,
12'hf86,
12'hf91,
12'hf94,
12'hf93,
12'hf9d,
12'hfbe,
12'h00e,
12'h077,
12'h0c1,
12'h0d2,
12'h0a2,
12'h060,
12'h042,
12'h068,
12'h0be,
12'h115,
12'h15a,
12'h164,
12'h13a,
12'h109,
12'h0ed,
12'h0ef,
12'h112,
12'h13c,
12'h146,
12'h12f,
12'h103,
12'h0d8,
12'h0b8,
12'h0a7,
12'h0a2,
12'h0b9,
12'h0de,
12'h0ea,
12'h0da,
12'h0b8,
12'h0b1,
12'h0be,
12'h0b9,
12'h096,
12'h05a,
12'h027,
12'h007,
12'hff5,
12'hff9,
12'h011,
12'h037,
12'h045,
12'h01a,
12'hfbf,
12'hf47,
12'hee7,
12'heb8,
12'heac,
12'hea9,
12'he9f,
12'he9d,
12'head,
12'hed0,
12'hef8,
12'hf0d,
12'hf17,
12'hf10,
12'hee8,
12'he9a,
12'he43,
12'he26,
12'he24,
12'he0a,
12'he02,
12'he32,
12'he89,
12'hed4,
12'hefa,
12'hf19,
12'hf55,
12'hf82,
12'hf53,
12'hed7,
12'he73,
12'he5f,
12'he71,
12'he62,
12'he38,
12'he27,
12'he46,
12'he95,
12'hef0,
12'hf4c,
12'hfa9,
12'hfdd,
12'hfc2,
12'hf64,
12'hf12,
12'hef8,
12'hef5,
12'hed9,
12'he9b,
12'he7f,
12'heb1,
12'hf0f,
12'hf7f,
12'hffa,
12'h077,
12'h0da,
12'h0ef,
12'h0b6,
12'h067,
12'h027,
12'hfee,
12'hfb4,
12'hf90,
12'hf99,
12'hfeb,
12'h08b,
12'h158,
12'h1fe,
12'h24a,
12'h256,
12'h23b,
12'h21b,
12'h1fa,
12'h1c7,
12'h1a4,
12'h1a0,
12'h1c1,
12'h1ee,
12'h213,
12'h26f,
12'h2f9,
12'h361,
12'h361,
12'h2fb,
12'h27a,
12'h209,
12'h1d1,
12'h1ec,
12'h22c,
12'h266,
12'h274,
12'h248,
12'h221,
12'h201,
12'h1d7,
12'h1b1,
12'h194,
12'h172,
12'h138,
12'h0fe,
12'h0d1,
12'h0a2,
12'h078,
12'h059,
12'h04d,
12'h058,
12'h069,
12'h082,
12'h09b,
12'h095,
12'h04a,
12'hfb0,
12'heec,
12'he3f,
12'he01,
12'he36,
12'hea3,
12'hf19,
12'hf71,
12'hfa7,
12'hfae,
12'hf91,
12'hf6a,
12'hf45,
12'hf11,
12'heac,
12'he34,
12'hdda,
12'hdc5,
12'hdfa,
12'he51,
12'heae,
12'heeb,
12'hef0,
12'hece,
12'hea6,
12'he98,
12'heac,
12'hecc,
12'hef6,
12'hf21,
12'hf2d,
12'hf16,
12'hef2,
12'hef9,
12'hf23,
12'hf40,
12'hf3d,
12'hf39,
12'hf4e,
12'hf70,
12'hfa6,
12'hfd5,
12'hfd6,
12'hfb1,
12'hf80,
12'hf5e,
12'hf50,
12'hf5e,
12'hf9b,
12'h001,
12'h068,
12'h08b,
12'h07e,
12'h087,
12'h0ab,
12'h0d0,
12'h0d7,
12'h0d8,
12'h0f2,
12'h114,
12'h12d,
12'h13a,
12'h14f,
12'h161,
12'h15c,
12'h14d,
12'h148,
12'h151,
12'h159,
12'h14d,
12'h136,
12'h119,
12'h0eb,
12'h0b5,
12'h09e,
12'h0aa,
12'h0cb,
12'h0ef,
12'h105,
12'h10d,
12'h109,
12'h0f5,
12'h0d1,
12'h0a3,
12'h06e,
12'h03c,
12'h00f,
12'hfec,
12'hfca,
12'hfc2,
12'hfe2,
12'h00a,
12'h02f,
12'h029,
12'hfea,
12'hf8f,
12'hf37,
12'hef7,
12'hecf,
12'heb3,
12'he8f,
12'he64,
12'he4c,
12'he68,
12'hea4,
12'hecd,
12'hec6,
12'he94,
12'he68,
12'he67,
12'he6f,
12'he66,
12'he53,
12'he51,
12'he5f,
12'he4f,
12'he3f,
12'he71,
12'hedc,
12'hf40,
12'hf77,
12'hf87,
12'hf75,
12'hf3d,
12'hed9,
12'he67,
12'he2f,
12'he45,
12'he7d,
12'he9e,
12'hea1,
12'heaf,
12'hee4,
12'hf2b,
12'hf5f,
12'hf77,
12'hf67,
12'hf29,
12'heca,
12'he90,
12'hea9,
12'hefa,
12'hf5c,
12'hf9c,
12'hfc0,
12'hff0,
12'h045,
12'h091,
12'h09e,
12'h070,
12'h026,
12'hfe2,
12'hfb9,
12'hfd6,
12'h02b,
12'h088,
12'h0b5,
12'h0c4,
12'h0e6,
12'h11a,
12'h156,
12'h188,
12'h1ad,
12'h1c6,
12'h1ae,
12'h166,
12'h13b,
12'h161,
12'h1cf,
12'h258,
12'h2ba,
12'h2ef,
12'h30b,
12'h306,
12'h2fb,
12'h2f8,
12'h2fd,
12'h2f9,
12'h2bc,
12'h258,
12'h1e5,
12'h185,
12'h178,
12'h1a8,
12'h1e5,
12'h1fe,
12'h1d1,
12'h178,
12'h125,
12'h109,
12'h124,
12'h14c,
12'h15c,
12'h131,
12'h0be,
12'h033,
12'hfdc,
12'hfe4,
12'h03b,
12'h092,
12'h08b,
12'h00a,
12'hf6a,
12'hf12,
12'hf1d,
12'hf6b,
12'hfb0,
12'hfa5,
12'hf36,
12'he95,
12'he0e,
12'he00,
12'he7a,
12'hf17,
12'hf80,
12'hf80,
12'hf25,
12'hea0,
12'he2e,
12'he19,
12'he67,
12'hec4,
12'hedc,
12'hea7,
12'he5b,
12'he35,
12'he49,
12'he88,
12'hede,
12'hf2e,
12'hf55,
12'hf39,
12'hee3,
12'heb1,
12'hecc,
12'hf02,
12'hf2b,
12'hf2f,
12'hf24,
12'hf19,
12'hf12,
12'hf2a,
12'hf81,
12'hffa,
12'h047,
12'h03a,
12'hfe1,
12'hf81,
12'hf4f,
12'hf59,
12'hf8f,
12'hfe5,
12'h032,
12'h03f,
12'h01b,
12'h00b,
12'h03e,
12'h08f,
12'h0d2,
12'h0ef,
12'h0ee,
12'h0ec,
12'h0e6,
12'h0e6,
12'h0fd,
12'h138,
12'h184,
12'h1ac,
12'h19c,
12'h158,
12'h105,
12'h0cf,
12'h0c4,
12'h0df,
12'h104,
12'h111,
12'h104,
12'h0ed,
12'h0c5,
12'h096,
12'h09f,
12'h0df,
12'h113,
12'h108,
12'h0c1,
12'h07e,
12'h05d,
12'h04d,
12'h048,
12'h051,
12'h068,
12'h061,
12'h02e,
12'hfed,
12'hfbf,
12'hfb5,
12'hfbc,
12'hfc8,
12'hfc5,
12'hf93,
12'hf21,
12'he9f,
12'he4c,
12'he36,
12'he50,
12'he78,
12'he89,
12'he87,
12'he74,
12'he4e,
12'he3a,
12'he54,
12'he9b,
12'hede,
12'hee5,
12'heab,
12'he64,
12'he44,
12'he40,
12'he5e,
12'he96,
12'hed8,
12'hf11,
12'hf26,
12'hf20,
12'hf20,
12'hf2f,
12'hf33,
12'hf0c,
12'hecb,
12'he95,
12'he85,
12'he8b,
12'he86,
12'he7d,
12'he99,
12'hef6,
12'hf65,
12'hfa8,
12'hfaa,
12'hf75,
12'hf1d,
12'hebf,
12'hea9,
12'heef,
12'hf62,
12'hfb7,
12'hfc0,
12'hfc2,
12'h000,
12'h071,
12'h0e9,
12'h127,
12'h108,
12'h082,
12'hfd6,
12'hf68,
12'hf68,
12'hfda,
12'h071,
12'h0d1,
12'h0ed,
12'h0f7,
12'h113,
12'h150,
12'h1a6,
12'h1fb,
12'h232,
12'h217,
12'h1ab,
12'h14d,
12'h159,
12'h1dc,
12'h281,
12'h2f1,
12'h327,
12'h32b,
12'h302,
12'h2cf,
12'h2a8,
12'h286,
12'h25b,
12'h215,
12'h1c4,
12'h18c,
12'h180,
12'h1a6,
12'h1d9,
12'h200,
12'h20b,
12'h1e9,
12'h1b5,
12'h190,
12'h170,
12'h141,
12'h0f4,
12'h09a,
12'h04f,
12'h022,
12'h019,
12'h024,
12'h042,
12'h065,
12'h06a,
12'h03c,
12'hff7,
12'hfc5,
12'hfa4,
12'hf6f,
12'hf10,
12'heb0,
12'he81,
12'he88,
12'heb7,
12'heff,
12'hf4e,
12'hf79,
12'hf5c,
12'hf11,
12'hed3,
12'heb9,
12'he9c,
12'he66,
12'he3d,
12'he33,
12'he34,
12'he36,
12'he64,
12'hec4,
12'hf14,
12'hf2f,
12'hf09,
12'hecd,
12'hec3,
12'hed7,
12'hef9,
12'hf19,
12'hf24,
12'hf18,
12'heee,
12'hec6,
12'hecc,
12'hf16,
12'hf7c,
12'hfc9,
12'hfe3,
12'hfc8,
12'hfad,
12'hfbc,
12'hfec,
12'h011,
12'h015,
12'hffb,
12'hfc1,
12'hf88,
12'hf83,
12'hfbd,
12'h025,
12'h089,
12'h0c4,
12'h0d5,
12'h0c9,
12'h0ad,
12'h09c,
12'h0bc,
12'h0fc,
12'h131,
12'h132,
12'h110,
12'h107,
12'h121,
12'h148,
12'h160,
12'h157,
12'h145,
12'h130,
12'h114,
12'h0f1,
12'h0c7,
12'h0ac,
12'h095,
12'h081,
12'h087,
12'h0b1,
12'h0f0,
12'h128,
12'h12a,
12'h0ec,
12'h098,
12'h06e,
12'h067,
12'h04d,
12'h019,
12'hfe9,
12'hfca,
12'hfa1,
12'hf7e,
12'hf88,
12'hfba,
12'hfe1,
12'hfdd,
12'hfc3,
12'hf90,
12'hf38,
12'hecc,
12'he7a,
12'he5e,
12'he58,
12'he4c,
12'he44,
12'he4e,
12'he64,
12'he6f,
12'he73,
12'he76,
12'he84,
12'he99,
12'he95,
12'he77,
12'he62,
12'he69,
12'he81,
12'he91,
12'he9a,
12'heb9,
12'hef1,
12'hf36,
12'hf6d,
12'hf7d,
12'hf62,
12'hf28,
12'hed8,
12'he82,
12'he45,
12'he39,
12'he54,
12'he7c,
12'hec5,
12'hf34,
12'hfaa,
12'hffc,
12'h011,
12'hff6,
12'hfba,
12'hf80,
12'hf53,
12'hf34,
12'hf2b,
12'hf36,
12'hf4f,
12'hf6f,
12'hfa2,
12'hff9,
12'h059,
12'h093,
12'h089,
12'h05a,
12'h02d,
12'hffc,
12'hfcf,
12'hfc1,
12'hff2,
12'h03e,
12'h06a,
12'h08a,
12'h0de,
12'h162,
12'h1d8,
12'h21b,
12'h230,
12'h23d,
12'h239,
12'h1fc,
12'h19e,
12'h179,
12'h1c8,
12'h253,
12'h29d,
12'h2ad,
12'h2ca,
12'h2f4,
12'h30c,
12'h2ef,
12'h2bd,
12'h29a,
12'h273,
12'h23e,
12'h21c,
12'h21f,
12'h236,
12'h238,
12'h219,
12'h1e6,
12'h18e,
12'h123,
12'h0c8,
12'h0bb,
12'h10b,
12'h165,
12'h183,
12'h157,
12'h0f6,
12'h08c,
12'h03d,
12'h01c,
12'h02f,
12'h042,
12'h00b,
12'hf8f,
12'hf1f,
12'hefd,
12'hf1e,
12'hf3b,
12'hf4a,
12'hf42,
12'hefb,
12'he80,
12'he2c,
12'he5b,
12'hef6,
12'hf90,
12'hfba,
12'hf64,
12'hecf,
12'he3c,
12'hdd8,
12'hdd6,
12'he4f,
12'heef,
12'hf31,
12'heec,
12'he7a,
12'he43,
12'he69,
12'heb4,
12'hef6,
12'hf16,
12'hef6,
12'hea6,
12'he68,
12'he85,
12'heff,
12'hf82,
12'hfb5,
12'hf84,
12'hf19,
12'hecc,
12'hedb,
12'hf4b,
12'hfe8,
12'h05e,
12'h078,
12'h02e,
12'hfa2,
12'hf32,
12'hf25,
12'hf59,
12'hfa5,
12'hfe4,
12'h00c,
12'h018,
12'h001,
12'h001,
12'h044,
12'h0b4,
12'h100,
12'h0f1,
12'h0a8,
12'h077,
12'h08d,
12'h0e1,
12'h14d,
12'h1a6,
12'h1c7,
12'h196,
12'h11a,
12'h09d,
12'h075,
12'h0ae,
12'h117,
12'h15f,
12'h161,
12'h12e,
12'h0e7,
12'h0b5,
12'h0a9,
12'h0c1,
12'h0eb,
12'h0fb,
12'h0e6,
12'h0c3,
12'h0a6,
12'h0a4,
12'h0a1,
12'h086,
12'h05e,
12'h03a,
12'h01a,
12'hff8,
12'hfd2,
12'hfb4,
12'hfbc,
12'hfd6,
12'hfe3,
12'hfc8,
12'hf8c,
12'hf3e,
12'hedf,
12'he8c,
12'he6e,
12'he8d,
12'heb8,
12'hebb,
12'he9d,
12'he82,
12'he7c,
12'he80,
12'he86,
12'he9d,
12'head,
12'he9e,
12'he6b,
12'he1d,
12'hdfd,
12'he1f,
12'he61,
12'hea4,
12'hee1,
12'hf20,
12'hf4e,
12'hf63,
12'hf65,
12'hf56,
12'hf29,
12'hee6,
12'he96,
12'he57,
12'he51,
12'he73,
12'hea0,
12'heba,
12'hed6,
12'hf1b,
12'hf8a,
12'hfe2,
12'hfe7,
12'hfa9,
12'hf48,
12'hedf,
12'hea3,
12'heaf,
12'hef0,
12'hf45,
12'hf72,
12'hf82,
12'hfb2,
12'h01d,
12'h0b5,
12'h121,
12'h12c,
12'h0c7,
12'h01f,
12'hf90,
12'hf5c,
12'hf8c,
12'hff9,
12'h06a,
12'h0bc,
12'h0f4,
12'h128,
12'h171,
12'h1d2,
12'h22e,
12'h26d,
12'h26a,
12'h20c,
12'h17c,
12'h119,
12'h133,
12'h1c2,
12'h275,
12'h2fd,
12'h33a,
12'h33c,
12'h31f,
12'h301,
12'h2e4,
12'h2bd,
12'h282,
12'h22e,
12'h1d7,
12'h19d,
12'h197,
12'h1d0,
12'h221,
12'h25c,
12'h26e,
12'h240,
12'h1e5,
12'h17c,
12'h123,
12'h0ee,
12'h0e5,
12'h0d6,
12'h09a,
12'h035,
12'hfdc,
12'hfd2,
12'h013,
12'h071,
12'h0a5,
12'h094,
12'h044,
12'hfd7,
12'hf7c,
12'hf37,
12'hf04,
12'hecb,
12'he87,
12'he55,
12'he47,
12'he6c,
12'hece,
12'hf45,
12'hf89,
12'hf85,
12'hf4f,
12'hefe,
12'heab,
12'he6a,
12'he49,
12'he44,
12'he44,
12'he44,
12'he5e,
12'he8e,
12'hec6,
12'heec,
12'hef1,
12'heee,
12'hef0,
12'hef1,
12'hedb,
12'hec9,
12'hee0,
12'hf0f,
12'hf1f,
12'hf0c,
12'hf10,
12'hf47,
12'hf7f,
12'hf95,
12'hf97,
12'hfa9,
12'hfc8,
12'hfe4,
12'hfed,
12'hfcf,
12'hfac,
12'hf92,
12'hf78,
12'hf60,
12'hf67,
12'hfa7,
12'hffd,
12'h050,
12'h096,
12'h0ba,
12'h0ca,
12'h0d0,
12'h0d1,
12'h0e4,
12'h0fe,
12'h10a,
12'h0fc,
12'h0e5,
12'h0f3,
12'h123,
12'h157,
12'h168,
12'h159,
12'h14d,
12'h138,
12'h114,
12'h0e4,
12'h0b7,
12'h09d,
12'h084,
12'h066,
12'h064,
12'h096,
12'h0e9,
12'h12c,
12'h13c,
12'h114,
12'h0d8,
12'h0a8,
12'h074,
12'h046,
12'h022,
12'hffe,
12'hfdb,
12'hfbc,
12'hfa3,
12'hf9e,
12'hfbf,
12'hff4,
12'h00f,
12'hffa,
12'hfac,
12'hf2d,
12'hea7,
12'he61,
12'he69,
12'he8a,
12'he99,
12'he8d,
12'he69,
12'he50,
12'he52,
12'he68,
12'he84,
12'he90,
12'hea6,
12'heb6,
12'he97,
12'he62,
12'he4f,
12'he76,
12'heac,
12'hed0,
12'hee6,
12'hf08,
12'hf35,
12'hf52,
12'hf5a,
12'hf5a,
12'hf59,
12'hf3d,
12'hedb,
12'he5c,
12'he05,
12'hdde,
12'hdf5,
12'he52,
12'hef0,
12'hf9b,
12'hffa,
12'hff8,
12'hfc4,
12'hf8c,
12'hf5e,
12'hf38,
12'hf1d,
12'hf0b,
12'hef1,
12'hed6,
12'heeb,
12'hf5b,
12'h00b,
12'h0a3,
12'h0e0,
12'h0b3,
12'h052,
12'hff0,
12'hfa8,
12'hfa6,
12'hfe0,
12'h028,
12'h056,
12'h050,
12'h043,
12'h087,
12'h11c,
12'h1a6,
12'h1ea,
12'h1e5,
12'h1c3,
12'h1b1,
12'h1a1,
12'h198,
12'h1bf,
12'h217,
12'h26b,
12'h280,
12'h271,
12'h290,
12'h2f4,
12'h353,
12'h355,
12'h303,
12'h28c,
12'h202,
12'h1ae,
12'h1bb,
12'h206,
12'h243,
12'h238,
12'h1fd,
12'h1c6,
12'h1a0,
12'h17f,
12'h169,
12'h16f,
12'h17f,
12'h159,
12'h0f0,
12'h07e,
12'h04b,
12'h050,
12'h06b,
12'h086,
12'h08b,
12'h060,
12'h000,
12'hfbc,
12'hfc0,
12'hfec,
12'hfea,
12'hf87,
12'hf05,
12'heb2,
12'he7f,
12'he60,
12'he7a,
12'hef4,
12'hf8d,
12'hfc2,
12'hf79,
12'hef8,
12'heaa,
12'he9c,
12'he96,
12'he94,
12'hea2,
12'heb2,
12'hea4,
12'he85,
12'he80,
12'he9b,
12'hec9,
12'heeb,
12'hef1,
12'hede,
12'hec5,
12'heb4,
12'hed3,
12'hf34,
12'hf95,
12'hfad,
12'hf65,
12'hf0d,
12'hedc,
12'hed5,
12'hf0e,
12'hf8e,
12'h00b,
12'h048,
12'h029,
12'hfc9,
12'hf6c,
12'hf4e,
12'hf87,
12'hfd2,
12'hfe7,
12'hfcb,
12'hfb5,
12'hfca,
12'h002,
12'h05d,
12'h0cd,
12'h11f,
12'h123,
12'h0c9,
12'h055,
12'h039,
12'h09f,
12'h144,
12'h1c4,
12'h1e8,
12'h1ae,
12'h133,
12'h0aa,
12'h06b,
12'h09f,
12'h122,
12'h181,
12'h174,
12'h117,
12'h0ad,
12'h075,
12'h07a,
12'h0c0,
12'h109,
12'h10d,
12'h0c6,
12'h05f,
12'h024,
12'h03a,
12'h085,
12'h0cc,
12'h0de,
12'h0a8,
12'h03e,
12'hfd0,
12'hf8f,
12'hf8f,
12'hfbc,
12'hfee,
12'hffe,
12'hfd4,
12'hf76,
12'hf22,
12'heed,
12'hecc,
12'hebd,
12'heb1,
12'he95,
12'he5b,
12'he2a,
12'he35,
12'he83,
12'hee4,
12'hf15,
12'hf07,
12'heca,
12'he87,
12'he5d,
12'he46,
12'he3a,
12'he3f,
12'he58,
12'he74,
12'he9e,
12'hee4,
12'hf3e,
12'hf89,
12'hfa7,
12'hf8e,
12'hf43,
12'hef7,
12'heb8,
12'he76,
12'he4f,
12'he51,
12'he5a,
12'he51,
12'he63,
12'hec0,
12'hf60,
12'hfe3,
12'h000,
12'hfd6,
12'hf80,
12'hf23,
12'hee8,
12'hee3,
12'hef7,
12'hefc,
12'heec,
12'hee3,
12'hf29,
12'hfc4,
12'h06b,
12'h0d7,
12'h0ea,
12'h0ab,
12'h03a,
12'hfd3,
12'hfae,
12'hfe2,
12'h022,
12'h03e,
12'h02d,
12'h022,
12'h071,
12'h10c,
12'h1a7,
12'h200,
12'h20e,
12'h1e0,
12'h18d,
12'h14d,
12'h156,
12'h1bf,
12'h25b,
12'h2c1,
12'h2d8,
12'h2c2,
12'h2b9,
12'h2ea,
12'h317,
12'h31f,
12'h2ea,
12'h274,
12'h1e9,
12'h191,
12'h194,
12'h1cc,
12'h219,
12'h255,
12'h25e,
12'h231,
12'h1f7,
12'h1c0,
12'h187,
12'h153,
12'h11f,
12'h0ea,
12'h0b0,
12'h076,
12'h031,
12'h001,
12'h00b,
12'h037,
12'h05f,
12'h07b,
12'h089,
12'h081,
12'h05b,
12'h009,
12'hf87,
12'hef0,
12'he7f,
12'he56,
12'he6a,
12'he96,
12'hec5,
12'hf09,
12'hf45,
12'hf69,
12'hf77,
12'hf64,
12'hf49,
12'hf1c,
12'hed4,
12'he85,
12'he4a,
12'he39,
12'he46,
12'he60,
12'he90,
12'hebc,
12'hecf,
12'hecd,
12'hecc,
12'hefd,
12'hf40,
12'hf59,
12'hf4d,
12'hf2c,
12'hf1a,
12'hf0c,
12'hef6,
12'hf09,
12'hf3c,
12'hf65,
12'hf6f,
12'hf62,
12'hf79,
12'hfbb,
12'h006,
12'h01d,
12'hfe5,
12'hfa1,
12'hf87,
12'hf8d,
12'hf9a,
12'hfb2,
12'hfe7,
12'h022,
12'h03f,
12'h055,
12'h06e,
12'h09b,
12'h0df,
12'h100,
12'h0ef,
12'h0d0,
12'h0d3,
12'h0f5,
12'h111,
12'h11a,
12'h117,
12'h11b,
12'h11c,
12'h124,
12'h148,
12'h176,
12'h187,
12'h161,
12'h0fd,
12'h088,
12'h03f,
12'h037,
12'h064,
12'h0a5,
12'h0d8,
12'h0ef,
12'h0e2,
12'h0d2,
12'h0cf,
12'h0d0,
12'h0b5,
12'h065,
12'h00c,
12'hfcf,
12'hfb5,
12'hfc4,
12'hfea,
12'h008,
12'h00d,
12'hffc,
12'hfcf,
12'hf91,
12'hf59,
12'hf2e,
12'hf0a,
12'hef4,
12'hee0,
12'hec2,
12'he9c,
12'he81,
12'he82,
12'he8e,
12'he9c,
12'hea1,
12'he97,
12'he94,
12'heac,
12'hed9,
12'heed,
12'hed3,
12'hea1,
12'he7f,
12'he80,
12'he90,
12'hea3,
12'heda,
12'hf2f,
12'hf75,
12'hf8a,
12'hf6c,
12'hf45,
12'hf27,
12'hef3,
12'hea4,
12'he42,
12'hde7,
12'hdc5,
12'he12,
12'hec8,
12'hf9d,
12'h027,
12'h043,
12'h000,
12'hf8c,
12'hf3e,
12'hf24,
12'hf1d,
12'hf10,
12'hee8,
12'hebd,
12'heba,
12'hf06,
12'hfa9,
12'h05e,
12'h0d9,
12'h0e6,
12'h099,
12'h034,
12'hfd4,
12'hf9e,
12'hfa9,
12'hfd0,
12'hffa,
12'h011,
12'h028,
12'h080,
12'h10b,
12'h18f,
12'h1e0,
12'h1f9,
12'h1f9,
12'h1f9,
12'h1e9,
12'h1b7,
12'h19e,
12'h1cf,
12'h231,
12'h26a,
12'h277,
12'h29a,
12'h2dc,
12'h318,
12'h324,
12'h2fe,
12'h2b7,
12'h261,
12'h218,
12'h1f7,
12'h1f5,
12'h1f8,
12'h1ec,
12'h1d3,
12'h1bc,
12'h19f,
12'h16e,
12'h13e,
12'h140,
12'h172,
12'h195,
12'h175,
12'h118,
12'h0a3,
12'h03a,
12'h012,
12'h034,
12'h06a,
12'h06d,
12'h01c,
12'hfae,
12'hf6b,
12'hf6a,
12'hf7b,
12'hf6c,
12'hf32,
12'hee2,
12'he8f,
12'he52,
12'he6e,
12'hf06,
12'hfbc,
12'hff7,
12'hf96,
12'hee8,
12'he52,
12'he13,
12'he1e,
12'he52,
12'he91,
12'hebc,
12'heb0,
12'he79,
12'he61,
12'he85,
12'hec2,
12'hee6,
12'heca,
12'he9b,
12'he8a,
12'he9a,
12'hec9,
12'hf17,
12'hf60,
12'hf66,
12'hf16,
12'heb9,
12'he90,
12'heb6,
12'hf3b,
12'hfdd,
12'h054,
12'h06c,
12'h01c,
12'hfa2,
12'hf40,
12'hf2a,
12'hf61,
12'hfaa,
12'hfc4,
12'hfb3,
12'hfb3,
12'hfe4,
12'h03a,
12'h09c,
12'h0f0,
12'h120,
12'h10c,
12'h0a4,
12'h039,
12'h03f,
12'h0c6,
12'h179,
12'h1ed,
12'h1f6,
12'h1a9,
12'h133,
12'h0cb,
12'h09d,
12'h0bb,
12'h104,
12'h13f,
12'h145,
12'h116,
12'h0e0,
12'h0c9,
12'h0de,
12'h104,
12'h102,
12'h0dd,
12'h0aa,
12'h087,
12'h087,
12'h096,
12'h0b0,
12'h0bc,
12'h0ad,
12'h08c,
12'h059,
12'h02e,
12'h004,
12'hfcc,
12'hfa0,
12'hfa0,
12'hfc3,
12'hfd5,
12'hfb8,
12'hf90,
12'hf5b,
12'hf0f,
12'hecd,
12'heac,
12'hea7,
12'he9b,
12'he7b,
12'he6e,
12'he93,
12'hed1,
12'hefb,
12'hefc,
12'heda,
12'heb2,
12'he90,
12'he5b,
12'he26,
12'he1b,
12'he2d,
12'he4c,
12'he77,
12'hecb,
12'hf47,
12'hf99,
12'hf98,
12'hf65,
12'hf29,
12'hefa,
12'hec6,
12'he83,
12'he56,
12'he58,
12'he64,
12'he6b,
12'he89,
12'hee8,
12'hf76,
12'hfcc,
12'hfb9,
12'hf76,
12'hf2f,
12'hef5,
12'hef1,
12'hf13,
12'hf36,
12'hf3d,
12'hf27,
12'hf22,
12'hf5f,
12'hfe1,
12'h06a,
12'h0bb,
12'h0b0,
12'h054,
12'hfec,
12'hf9e,
12'hfa4,
12'hff1,
12'h03c,
12'h062,
12'h054,
12'h04e,
12'h082,
12'h0fc,
12'h1a4,
12'h224,
12'h242,
12'h1f2,
12'h170,
12'h11a,
12'h112,
12'h166,
12'h1fc,
12'h28e,
12'h2e6,
12'h301,
12'h308,
12'h315,
12'h31c,
12'h313,
12'h2dc,
12'h26d,
12'h1f7,
12'h19b,
12'h17b,
12'h19e,
12'h1eb,
12'h241,
12'h25b,
12'h22c,
12'h1d7,
12'h190,
12'h16a,
12'h158,
12'h164,
12'h168,
12'h141,
12'h0f1,
12'h082,
12'h044,
12'h04c,
12'h060,
12'h058,
12'h01e,
12'hfd7,
12'hfae,
12'hfc2,
12'hffb,
12'h014,
12'hfeb,
12'hf74,
12'hedb,
12'he59,
12'he12,
12'he2d,
12'hea3,
12'hf23,
12'hf65,
12'hf4f,
12'hf13,
12'heeb,
12'hedb,
12'hedb,
12'hecb,
12'hea1,
12'he76,
12'he58,
12'he51,
12'he67,
12'he9c,
12'hedb,
12'hefd,
12'hefa,
12'heda,
12'heaf,
12'he89,
12'he90,
12'hece,
12'hf1d,
12'hf4e,
12'hf46,
12'hf2c,
12'hf2d,
12'hf4c,
12'hf7a,
12'hfa7,
12'hfd2,
12'hfe8,
12'hfdd,
12'hfbb,
12'hf96,
12'hf98,
12'hfca,
12'h000,
12'h00e,
12'hffb,
12'hfdb,
12'hfd0,
12'hfff,
12'h053,
12'h0b7,
12'h105,
12'h116,
12'h0ea,
12'h0a9,
12'h090,
12'h0c8,
12'h134,
12'h180,
12'h181,
12'h13f,
12'h0e6,
12'h0b4,
12'h0c7,
12'h11a,
12'h173,
12'h192,
12'h15a,
12'h0e8,
12'h07a,
12'h03e,
12'h041,
12'h06e,
12'h0a4,
12'h0c2,
12'h0b1,
12'h082,
12'h069,
12'h08d,
12'h0c3,
12'h0c9,
12'h08b,
12'h029,
12'hfbd,
12'hf64,
12'hf47,
12'hf5d,
12'hfa6,
12'hffc,
12'h025,
12'h007,
12'hfab,
12'hf4d,
12'hefb,
12'hec9,
12'hebe,
12'heb5,
12'heb1,
12'hea5,
12'he88,
12'he71,
12'he71,
12'he89,
12'hea2,
12'hea2,
12'he97,
12'he99,
12'he9c,
12'he8c,
12'he6d,
12'he5e,
12'he75,
12'he9d,
12'hec0,
12'hee8,
12'hf1d,
12'hf4d,
12'hf51,
12'hf30,
12'hf0e,
12'hefa,
12'hefd,
12'hee9,
12'heab,
12'he5d,
12'he21,
12'he18,
12'he55,
12'hee8,
12'hf8e,
12'hff0,
12'hff5,
12'hfb4,
12'hf70,
12'hf54,
12'hf63,
12'hf72,
12'hf5a,
12'hf1b,
12'hed6,
12'hecf,
12'hf31,
12'hfd1,
12'h062,
12'h09b,
12'h06f,
12'h013,
12'hfc1,
12'hfae,
12'hfd4,
12'h00d,
12'h03f,
12'h04f,
12'h03e,
12'h039,
12'h07b,
12'h0fd,
12'h177,
12'h1b3,
12'h1b2,
12'h19d,
12'h19c,
12'h1b1,
12'h1d4,
12'h218,
12'h279,
12'h2bb,
12'h2c0,
12'h2b3,
12'h2be,
12'h2df,
12'h302,
12'h2fe,
12'h2c0,
12'h259,
12'h1fc,
12'h1d9,
12'h1fa,
12'h238,
12'h251,
12'h23f,
12'h226,
12'h205,
12'h1db,
12'h1a1,
12'h177,
12'h175,
12'h175,
12'h15e,
12'h124,
12'h0d9,
12'h097,
12'h077,
12'h07b,
12'h08d,
12'h08c,
12'h058,
12'h010,
12'hfef,
12'hff4,
12'hfe7,
12'hf9d,
12'hf2c,
12'hec5,
12'he76,
12'he4a,
12'he51,
12'heb1,
12'hf56,
12'hfc6,
12'hfbe,
12'hf57,
12'hed6,
12'he82,
12'he71,
12'he82,
12'he98,
12'hea8,
12'hea3,
12'he7c,
12'he52,
12'he58,
12'he8a,
12'hec1,
12'hecf,
12'heb0,
12'he7e,
12'he56,
12'he60,
12'heb6,
12'hf42,
12'hfb0,
12'hfa8,
12'hf4b,
12'heee,
12'hece,
12'hef8,
12'hf4e,
12'hfb1,
12'hfed,
12'hfe6,
12'hfab,
12'hf70,
12'hf67,
12'hfa1,
12'hfff,
12'h025,
12'hfec,
12'hf93,
12'hf66,
12'hf91,
12'h002,
12'h083,
12'h0ed,
12'h114,
12'h0e8,
12'h088,
12'h047,
12'h076,
12'h106,
12'h1a1,
12'h1ee,
12'h1c3,
12'h148,
12'h0d2,
12'h0b8,
12'h0fc,
12'h16a,
12'h1af,
12'h19f,
12'h14a,
12'h0d9,
12'h094,
12'h08e,
12'h0be,
12'h106,
12'h121,
12'h0fa,
12'h0ac,
12'h06f,
12'h06e,
12'h0a4,
12'h0dd,
12'h0e5,
12'h0a1,
12'h03c,
12'hff3,
12'hfd4,
12'hfd7,
12'hfdd,
12'hfe2,
12'hfec,
12'hfe7,
12'hfc2,
12'hf7d,
12'hf31,
12'hef8,
12'hed9,
12'hed8,
12'hedf,
12'hec5,
12'he99,
12'he81,
12'he7f,
12'he8c,
12'he99,
12'he9d,
12'he9d,
12'he86,
12'he6a,
12'he65,
12'he64,
12'he4b,
12'he20,
12'he1e,
12'he5f,
12'hebb,
12'hef8,
12'hf15,
12'hf35,
12'hf58,
12'hf54,
12'hf20,
12'hef6,
12'hef3,
12'hee3,
12'he9d,
12'he42,
12'he0f,
12'he1e,
12'he5a,
12'hec3,
12'hf48,
12'hfaa,
12'hfce,
12'hfb4,
12'hf7a,
12'hf51,
12'hf38,
12'hf25,
12'hf07,
12'hecd,
12'he95,
12'he90,
12'hee1,
12'hf80,
12'h03a,
12'h0d4,
12'h107,
12'h0da,
12'h082,
12'h02b,
12'hff7,
12'hfe4,
12'hfe2,
12'hfea,
12'hff5,
12'h008,
12'h054,
12'h0f7,
12'h1bd,
12'h23b,
12'h23a,
12'h1ec,
12'h1a7,
12'h19a,
12'h1ae,
12'h1bd,
12'h1d9,
12'h216,
12'h24c,
12'h277,
12'h2b5,
12'h319,
12'h387,
12'h3ad,
12'h364,
12'h2d3,
12'h235,
12'h1c7,
12'h1c3,
12'h1f9,
12'h223,
12'h22d,
12'h212,
12'h1ef,
12'h1e3,
12'h1e8,
12'h1e1,
12'h1c6,
12'h190,
12'h138,
12'h0dc,
12'h0a1,
12'h095,
12'h09b,
12'h09b,
12'h07c,
12'h03d,
12'h016,
12'h01a,
12'h03d,
12'h055,
12'h038,
12'hfdf,
12'hf47,
12'he9c,
12'he3d,
12'he4d,
12'he98,
12'hee5,
12'hf16,
12'hf23,
12'hf1c,
12'hf07,
12'hf00,
12'hf2c,
12'hf69,
12'hf4e,
12'hebb,
12'he09,
12'hda3,
12'hda8,
12'hded,
12'he49,
12'hea4,
12'hee2,
12'hedc,
12'he97,
12'he75,
12'heaf,
12'hf0d,
12'hf41,
12'hf33,
12'hf02,
12'heca,
12'he91,
12'he7a,
12'hebe,
12'hf3d,
12'hf9c,
12'hfa3,
12'hf71,
12'hf4f,
12'hf68,
12'hfac,
12'hfd8,
12'hfe2,
12'hfde,
12'hfc4,
12'hf8c,
12'hf51,
12'hf60,
12'hfca,
12'h04c,
12'h09d,
12'h0a8,
12'h0a0,
12'h096,
12'h07a,
12'h060,
12'h075,
12'h0dc,
12'h15c,
12'h193,
12'h16f,
12'h126,
12'h0fe,
12'h0fe,
12'h114,
12'h141,
12'h17c,
12'h1a2,
12'h182,
12'h11c,
12'h0be,
12'h0a1,
12'h0b3,
12'h0db,
12'h0f8,
12'h0f2,
12'h0d4,
12'h0b0,
12'h0a2,
12'h0c3,
12'h0fa,
12'h113,
12'h0ea,
12'h080,
12'h002,
12'hfae,
12'hf92,
12'hfac,
12'hfe4,
12'h01d,
12'h027,
12'hfe9,
12'hf8c,
12'hf53,
12'hf56,
12'hf5a,
12'hf42,
12'hf1a,
12'hede,
12'hea2,
12'he61,
12'he3c,
12'he57,
12'he94,
12'hec8,
12'hec0,
12'he89,
12'he6f,
12'he87,
12'heb6,
12'hecd,
12'hebe,
12'hea2,
12'he8d,
12'he83,
12'he81,
12'hea5,
12'hefc,
12'hf5b,
12'hf82,
12'hf62,
12'hf2e,
12'hf0e,
12'hef9,
12'hed3,
12'he91,
12'he4e,
12'he25,
12'he29,
12'he79,
12'hf17,
12'hfc5,
12'h030,
12'h03c,
12'h00b,
12'hfdb,
12'hfbe,
12'hf8a,
12'hf2b,
12'hec5,
12'he87,
12'he86,
12'hebc,
12'hf27,
12'hfb7,
12'h045,
12'h0ad,
12'h0d3,
12'h0cb,
12'h0a4,
12'h057,
12'hff6,
12'hfac,
12'hf96,
12'hfb2,
12'hfea,
12'h032,
12'h0ac,
12'h150,
12'h1e0,
12'h22c,
12'h23e,
12'h24b,
12'h267,
12'h260,
12'h210,
12'h1b0,
12'h191,
12'h1c7,
12'h21d,
12'h26f,
12'h2d1,
12'h32b,
12'h34e,
12'h331,
12'h2ea,
12'h2a9,
12'h273,
12'h24e,
12'h236,
12'h20b,
12'h1d4,
12'h1a3,
12'h19e,
12'h1b6,
12'h1b8,
12'h1a4,
12'h198,
12'h19e,
12'h19b,
12'h178,
12'h146,
12'h112,
12'h0cc,
12'h072,
12'h01f,
12'hfeb,
12'hfe5,
12'hffa,
12'h01c,
12'h02c,
12'hffb,
12'hf99,
12'hf21,
12'heb4,
12'he72,
12'he66,
12'he8d,
12'hecb,
12'hf02,
12'hf33,
12'hf5e,
12'hf5e,
12'hf34,
12'hf0f,
12'hf06,
12'hee2,
12'he85,
12'he21,
12'he00,
12'he39,
12'he7c,
12'he89,
12'he8c,
12'he9e,
12'hea3,
12'he7b,
12'he38,
12'he32,
12'he84,
12'hef1,
12'hf34,
12'hf43,
12'hf2a,
12'hef7,
12'heb0,
12'he81,
12'he9b,
12'hee8,
12'hf38,
12'hf69,
12'hf84,
12'hf99,
12'hfa8,
12'hfb1,
12'hfab,
12'hf97,
12'hf84,
12'hf5a,
12'hf1b,
12'hf0a,
12'hf55,
12'hfde,
12'h04a,
12'h073,
12'h07c,
12'h08f,
12'h08b,
12'h053,
12'h03a,
12'h096,
12'h138,
12'h1a8,
12'h19d,
12'h13f,
12'h0fc,
12'h0ef,
12'h0f3,
12'h0fe,
12'h11a,
12'h135,
12'h13e,
12'h126,
12'h10a,
12'h119,
12'h136,
12'h144,
12'h131,
12'h0fc,
12'h0c5,
12'h0aa,
12'h0bb,
12'h0d8,
12'h0e2,
12'h0d6,
12'h0bb,
12'h08c,
12'h057,
12'h040,
12'h044,
12'h03c,
12'h00c,
12'hfd8,
12'hfc0,
12'hfbd,
12'hfa4,
12'hf80,
12'hf80,
12'hf90,
12'hf76,
12'hf21,
12'hecb,
12'he9e,
12'he8d,
12'he6f,
12'he5a,
12'he7e,
12'hecb,
12'hef4,
12'hed8,
12'hea2,
12'he81,
12'he7a,
12'he5c,
12'he2b,
12'he2f,
12'he7c,
12'hec6,
12'heda,
12'hedb,
12'hefc,
12'hf2a,
12'hf28,
12'hef8,
12'hece,
12'hecc,
12'hec9,
12'he95,
12'he51,
12'he3a,
12'he65,
12'hea2,
12'hedd,
12'hf3a,
12'hfa7,
12'hfe3,
12'hfcf,
12'hf92,
12'hf71,
12'hf75,
12'hf6c,
12'hf3b,
12'hef6,
12'hec8,
12'hece,
12'hf0c,
12'hf61,
12'hfcc,
12'h04d,
12'h0b0,
12'h0b7,
12'h062,
12'hff9,
12'hfa6,
12'hf82,
12'hf9a,
12'hfec,
12'h054,
12'h08d,
12'h097,
12'h0ca,
12'h163,
12'h22c,
12'h2b3,
12'h2b1,
12'h24c,
12'h1cd,
12'h15b,
12'h109,
12'h10a,
12'h191,
12'h254,
12'h2cc,
12'h2d3,
12'h2cd,
12'h313,
12'h371,
12'h38e,
12'h34d,
12'h2cd,
12'h235,
12'h1af,
12'h16e,
12'h18b,
12'h1d8,
12'h20e,
12'h218,
12'h1f8,
12'h1b8,
12'h18c,
12'h195,
12'h1bd,
12'h1d8,
12'h1b9,
12'h14c,
12'h0b3,
12'h029,
12'hff1,
12'h00b,
12'h03e,
12'h054,
12'h050,
12'h03c,
12'h009,
12'hfcf,
12'hfb9,
12'hfb8,
12'hf8c,
12'hf28,
12'hec7,
12'he8f,
12'he82,
12'he8d,
12'heb1,
12'hef4,
12'hf24,
12'hf2c,
12'hf22,
12'hf28,
12'hf39,
12'hf12,
12'heb9,
12'he72,
12'he61,
12'he72,
12'he71,
12'he74,
12'he99,
12'hebe,
12'heb8,
12'he8b,
12'he93,
12'heed,
12'hf43,
12'hf54,
12'hf2b,
12'heec,
12'heb5,
12'hea0,
12'hec2,
12'hf19,
12'hf6c,
12'hf87,
12'hf64,
12'hf38,
12'hf3d,
12'hf78,
12'hfb9,
12'hfcf,
12'hfb7,
12'hf8a,
12'hf55,
12'hf2f,
12'hf3c,
12'hf8b,
12'h009,
12'h05d,
12'h061,
12'h05b,
12'h073,
12'h0a2,
12'h0cc,
12'h0e9,
12'h115,
12'h138,
12'h12d,
12'h0f7,
12'h0c1,
12'h0bf,
12'h0eb,
12'h112,
12'h124,
12'h133,
12'h145,
12'h145,
12'h12f,
12'h10c,
12'h0da,
12'h0a7,
12'h079,
12'h065,
12'h080,
12'h0c4,
12'h110,
12'h13e,
12'h136,
12'h0f5,
12'h0a5,
12'h06f,
12'h05c,
12'h04a,
12'h02f,
12'h00a,
12'hfda,
12'hfb5,
12'hfbb,
12'hfdf,
12'hfef,
12'hfd2,
12'hf86,
12'hf37,
12'heff,
12'hef2,
12'hf0a,
12'hf1c,
12'hf0e,
12'hed2,
12'he85,
12'he52,
12'he54,
12'he85,
12'heb4,
12'heb4,
12'he8f,
12'he77,
12'he7c,
12'he7f,
12'he7a,
12'he91,
12'hec6,
12'hee6,
12'hed4,
12'heb6,
12'hebd,
12'hef8,
12'hf3f,
12'hf59,
12'hf3f,
12'hf0a,
12'hedd,
12'heae,
12'he77,
12'he5a,
12'he67,
12'he86,
12'heb7,
12'hf13,
12'hf8a,
12'hff2,
12'h022,
12'h00f,
12'hfc6,
12'hf73,
12'hf31,
12'hf12,
12'hf14,
12'hf17,
12'hf1c,
12'hf3c,
12'hf78,
12'hfbf,
12'h01d,
12'h08a,
12'h0cb,
12'h0ad,
12'h03f,
12'hfcf,
12'hf8a,
12'hf84,
12'hfc0,
12'h01f,
12'h07e,
12'h0b1,
12'h0cd,
12'h112,
12'h197,
12'h222,
12'h264,
12'h248,
12'h1fa,
12'h1a6,
12'h152,
12'h122,
12'h15c,
12'h1fa,
12'h282,
12'h2ad,
12'h2aa,
12'h2cb,
12'h31a,
12'h346,
12'h323,
12'h2d1,
12'h25a,
12'h1d9,
12'h182,
12'h176,
12'h1a4,
12'h1c3,
12'h1c2,
12'h1b0,
12'h190,
12'h179,
12'h174,
12'h17d,
12'h18b,
12'h174,
12'h118,
12'h08b,
12'h00f,
12'hfde,
12'hff6,
12'h02d,
12'h057,
12'h059,
12'h02e,
12'hff1,
12'hfc6,
12'hfc3,
12'hfc1,
12'hf86,
12'hf16,
12'hea6,
12'he68,
12'he52,
12'he73,
12'hee1,
12'hf59,
12'hf8a,
12'hf5d,
12'hf0b,
12'hedf,
12'hedc,
12'hecd,
12'hea3,
12'he83,
12'he87,
12'he9f,
12'hea3,
12'he9c,
12'heae,
12'hecb,
12'hecb,
12'heaf,
12'hea4,
12'hece,
12'hf0d,
12'hf34,
12'hf4c,
12'hf55,
12'hf2f,
12'hedd,
12'heaa,
12'hec6,
12'hf23,
12'hf80,
12'hfad,
12'hfc4,
12'hfbf,
12'hfae,
12'hfac,
12'hfaf,
12'hfbd,
12'hfd1,
12'hfca,
12'hf9a,
12'hf6a,
12'hf7f,
12'hfec,
12'h06a,
12'h0b0,
12'h0b7,
12'h0a8,
12'h0a7,
12'h0a2,
12'h09a,
12'h0cd,
12'h13b,
12'h193,
12'h195,
12'h14e,
12'h107,
12'h0ed,
12'h0e9,
12'h0e1,
12'h0fb,
12'h13b,
12'h16c,
12'h15b,
12'h10f,
12'h0c5,
12'h09d,
12'h089,
12'h082,
12'h099,
12'h0c5,
12'h0da,
12'h0d1,
12'h0be,
12'h0aa,
12'h099,
12'h093,
12'h08b,
12'h068,
12'h032,
12'hff7,
12'hfb9,
12'hf97,
12'hfa9,
12'hfda,
12'h005,
12'hff8,
12'hfb4,
12'hf74,
12'hf47,
12'hf20,
12'hf03,
12'heef,
12'hed1,
12'hea5,
12'he75,
12'he5e,
12'he76,
12'heb3,
12'hedd,
12'hecc,
12'hea2,
12'he8b,
12'he8f,
12'he85,
12'he67,
12'he56,
12'he69,
12'he92,
12'hea6,
12'hea4,
12'heca,
12'hf15,
12'hf4d,
12'hf68,
12'hf65,
12'hf54,
12'hf3c,
12'heec,
12'he75,
12'he3a,
12'he5f,
12'heac,
12'hec9,
12'hebe,
12'hee0,
12'hf40,
12'hf9b,
12'hfb6,
12'hfa7,
12'hf83,
12'hf2a,
12'hecb,
12'head,
12'hee3,
12'hf4e,
12'hf90,
12'hf9d,
12'hfbd,
12'h011,
12'h07d,
12'h0be,
12'h0ac,
12'h063,
12'h003,
12'hfad,
12'hf8e,
12'hfc8,
12'h049,
12'h0bb,
12'h0e9,
12'h0fa,
12'h10e,
12'h13a,
12'h17e,
12'h1c5,
12'h1f0,
12'h1d8,
12'h17a,
12'h10b,
12'h0ee,
12'h147,
12'h1f9,
12'h2ab,
12'h301,
12'h2ff,
12'h2e3,
12'h2d8,
12'h2e4,
12'h2f9,
12'h2e6,
12'h293,
12'h21c,
12'h1a0,
12'h13c,
12'h12a,
12'h17a,
12'h1ed,
12'h22f,
12'h210,
12'h1c0,
12'h18c,
12'h18c,
12'h19b,
12'h191,
12'h15c,
12'h0f6,
12'h069,
12'hfe9,
12'hfc6,
12'h008,
12'h07b,
12'h0b9,
12'h084,
12'h01c,
12'hfbe,
12'hf9f,
12'hfcb,
12'hfdd,
12'hfac,
12'hf49,
12'heb4,
12'he41,
12'he34,
12'he95,
12'hf2d,
12'hf91,
12'hf88,
12'hf21,
12'heb6,
12'he86,
12'he8b,
12'hea3,
12'hea7,
12'he9e,
12'he7f,
12'he51,
12'he32,
12'he5c,
12'hebe,
12'hf05,
12'hf06,
12'hed8,
12'hec1,
12'hec2,
12'hed7,
12'hefb,
12'hf22,
12'hf3d,
12'hf0c,
12'hea6,
12'he78,
12'hec2,
12'hf59,
12'hfd8,
12'h000,
12'hfdf,
12'hfb4,
12'hf93,
12'hf88,
12'hfa6,
12'hfd2,
12'hff1,
12'hfe0,
12'hfa5,
12'hf7d,
12'hf97,
12'hffa,
12'h087,
12'h0fe,
12'h128,
12'h103,
12'h0a8,
12'h06b,
12'h086,
12'h0de,
12'h14b,
12'h186,
12'h16e,
12'h12a,
12'h0f2,
12'h0ea,
12'h109,
12'h135,
12'h161,
12'h183,
12'h175,
12'h136,
12'h0ee,
12'h0bc,
12'h0a4,
12'h08f,
12'h07c,
12'h082,
12'h0ad,
12'h0dd,
12'h0f2,
12'h0df,
12'h0d6,
12'h0e8,
12'h0db,
12'h0a1,
12'h052,
12'h006,
12'hfc8,
12'hf89,
12'hf73,
12'hfa0,
12'hfe9,
12'h020,
12'h01f,
12'hfef,
12'hf9b,
12'hf22,
12'hea0,
12'he5f,
12'he7c,
12'hea6,
12'hea4,
12'he8a,
12'he76,
12'he76,
12'he8a,
12'he9f,
12'heba,
12'hed6,
12'hec6,
12'he90,
12'he53,
12'he43,
12'he74,
12'hea5,
12'hec7,
12'hecf,
12'hec4,
12'hebb,
12'heca,
12'hf09,
12'hf5a,
12'hf86,
12'hf6e,
12'hf16,
12'hea9,
12'he6b,
12'he6c,
12'he7c,
12'he7c,
12'he69,
12'he7d,
12'hee1,
12'hf5b,
12'hfb0,
12'hfb7,
12'hf8a,
12'hf45,
12'hef7,
12'hedf,
12'hf06,
12'hf54,
12'hf80,
12'hf6e,
12'hf77,
12'hfde,
12'h06f,
12'h0c5,
12'h0b1,
12'h060,
12'h00c,
12'hfb8,
12'hf87,
12'hfa2,
12'hffb,
12'h04f,
12'h06b,
12'h086,
12'h0db,
12'h151,
12'h1ad,
12'h1d4,
12'h1e0,
12'h1da,
12'h1a8,
12'h160,
12'h13f,
12'h18e,
12'h239,
12'h2ca,
12'h308,
12'h305,
12'h2e6,
12'h2cf,
12'h2cb,
12'h2c5,
12'h2a4,
12'h259,
12'h1ff,
12'h1be,
12'h1a6,
12'h1be,
12'h1e7,
12'h200,
12'h202,
12'h1d0,
12'h186,
12'h155,
12'h13e,
12'h137,
12'h12d,
12'h113,
12'h0f4,
12'h0c0,
12'h07e,
12'h04f,
12'h03b,
12'h046,
12'h058,
12'h05d,
12'h03e,
12'h006,
12'hfde,
12'hfb2,
12'hf6a,
12'hf1d,
12'hee6,
12'hec3,
12'hec5,
12'hedc,
12'hef8,
12'hf25,
12'hf4d,
12'hf59,
12'hf4a,
12'hf38,
12'hf28,
12'hee7,
12'he80,
12'he32,
12'he1b,
12'he37,
12'he68,
12'heb1,
12'heff,
12'hf15,
12'hed4,
12'he66,
12'he3a,
12'he77,
12'hed7,
12'hf0e,
12'hf1a,
12'hf0d,
12'hee2,
12'heaa,
12'he9d,
12'hef6,
12'hf7a,
12'hfbf,
12'hf9c,
12'hf3f,
12'hf1a,
12'hf5e,
12'hfda,
12'h043,
12'h05d,
12'h014,
12'hf85,
12'hefa,
12'hec8,
12'hf0e,
12'hfae,
12'h054,
12'h0bd,
12'h0cb,
12'h096,
12'h06a,
12'h073,
12'h0b8,
12'h116,
12'h156,
12'h14e,
12'h109,
12'h0c6,
12'h0c6,
12'h106,
12'h156,
12'h181,
12'h16f,
12'h140,
12'h109,
12'h0c9,
12'h098,
12'h08e,
12'h0a1,
12'h0a8,
12'h095,
12'h089,
12'h0a1,
12'h0d4,
12'h0fe,
12'h0f8,
12'h0cd,
12'h0b0,
12'h0a5,
12'h082,
12'h040,
12'h003,
12'hfef,
12'hff0,
12'hfed,
12'hfe5,
12'hfd4,
12'hfc8,
12'hfb8,
12'hfac,
12'hfab,
12'hf95,
12'hf53,
12'heec,
12'he9c,
12'he93,
12'hea5,
12'hea6,
12'he95,
12'he86,
12'he8a,
12'he98,
12'he9a,
12'heaa,
12'heca,
12'heda,
12'hebc,
12'he7d,
12'he50,
12'he4c,
12'he63,
12'he81,
12'hea2,
12'heca,
12'hf0d,
12'hf51,
12'hf70,
12'hf65,
12'hf35,
12'hf0b,
12'hee7,
12'hea7,
12'he61,
12'he31,
12'he34,
12'he7d,
12'hf01,
12'hf9a,
12'h002,
12'h022,
12'hffc,
12'hfb2,
12'hf7e,
12'hf72,
12'hf5c,
12'hf1a,
12'hebf,
12'he84,
12'hea2,
12'hf02,
12'hf91,
12'h033,
12'h0b7,
12'h0f0,
12'h0cd,
12'h0a0,
12'h09c,
12'h096,
12'h06a,
12'h00b,
12'hfb7,
12'hfa2,
12'hfc8,
12'h043,
12'h113,
12'h1f9,
12'h27d,
12'h265,
12'h213,
12'h200,
12'h217,
12'h20f,
12'h1df,
12'h1b6,
12'h1bd,
12'h1c8,
12'h1d1,
12'h218,
12'h2a8,
12'h32b,
12'h33d,
12'h2e3,
12'h26d,
12'h202,
12'h1c2,
12'h1dd,
12'h233,
12'h25b,
12'h21c,
12'h19a,
12'h142,
12'h150,
12'h17a,
12'h195,
12'h19b,
12'h184,
12'h132,
12'h0bc,
12'h080,
12'h093,
12'h0c9,
12'h0cf,
12'h082,
12'h010,
12'hfbf,
12'hfae,
12'hfc9,
12'hff0,
12'h00d,
12'hfe3,
12'hf57,
12'heb8,
12'he67,
12'he86,
12'hede,
12'hf30,
12'hf61,
12'hf74,
12'hf60,
12'hf2b,
12'hef2,
12'hee6,
12'hef1,
12'hec1,
12'he58,
12'hdfe,
12'hdf2,
12'he33,
12'he77,
12'he9d,
12'heba,
12'hed2,
12'hecb,
12'hea7,
12'hea2,
12'hed8,
12'hf20,
12'hf46,
12'hf40,
12'hf24,
12'hefb,
12'hecd,
12'he9d,
12'hea4,
12'hefd,
12'hf65,
12'hfa8,
12'hfb7,
12'hfae,
12'hfa9,
12'hf9d,
12'hf85,
12'hf69,
12'hf68,
12'hf7c,
12'hf7c,
12'hf7c,
12'hfb2,
12'h018,
12'h05f,
12'h064,
12'h05f,
12'h08b,
12'h0c8,
12'h0d5,
12'h0b4,
12'h0b5,
12'h104,
12'h15d,
12'h180,
12'h170,
12'h151,
12'h122,
12'h0d3,
12'h0a4,
12'h0c3,
12'h121,
12'h17b,
12'h184,
12'h140,
12'h0d7,
12'h084,
12'h079,
12'h0ab,
12'h0ef,
12'h108,
12'h0ec,
12'h0c1,
12'h0a7,
12'h0a6,
12'h0bd,
12'h0dd,
12'h0df,
12'h0a4,
12'h037,
12'hfe2,
12'hfd3,
12'hff6,
12'h028,
12'h03d,
12'h020,
12'hfce,
12'hf69,
12'hf3b,
12'hf48,
12'hf6c,
12'hf63,
12'hf14,
12'heb9,
12'he74,
12'he45,
12'he41,
12'he87,
12'hefe,
12'hf49,
12'hf21,
12'hea3,
12'he3c,
12'he24,
12'he49,
12'he63,
12'he66,
12'he78,
12'he8d,
12'he8b,
12'he8b,
12'hebf,
12'hf29,
12'hf8e,
12'hfb3,
12'hf8f,
12'hf32,
12'hece,
12'he87,
12'he5c,
12'he5c,
12'he95,
12'hec6,
12'heb2,
12'he72,
12'he6e,
12'hed8,
12'hf6f,
12'hfc4,
12'hfa7,
12'hf48,
12'hed9,
12'he7d,
12'he69,
12'heb3,
12'hf31,
12'hf8e,
12'hf97,
12'hf94,
12'hfd5,
12'h05c,
12'h0e6,
12'h105,
12'h0ae,
12'h013,
12'hf78,
12'hf1c,
12'hf25,
12'hf8e,
12'h012,
12'h06b,
12'h098,
12'h0cc,
12'h123,
12'h191,
12'h1f4,
12'h226,
12'h1fb,
12'h17b,
12'h0d5,
12'h072,
12'h0b5,
12'h18f,
12'h286,
12'h31f,
12'h33f,
12'h319,
12'h2fa,
12'h309,
12'h32c,
12'h32a,
12'h2e3,
12'h252,
12'h1a8,
12'h123,
12'h10b,
12'h166,
12'h1ef,
12'h258,
12'h244,
12'h1d1,
12'h171,
12'h166,
12'h195,
12'h1ca,
12'h1d5,
12'h197,
12'h0ed,
12'h00f,
12'hf86,
12'hfa7,
12'h044,
12'h0c4,
12'h0cd,
12'h065,
12'hfd5,
12'hf93,
12'hfd5,
12'h048,
12'h077,
12'h01d,
12'hf50,
12'he67,
12'hdda,
12'hdfe,
12'heba,
12'hf8c,
12'hfe8,
12'hfa2,
12'hefc,
12'he80,
12'he6b,
12'he9e,
12'hee2,
12'hf0c,
12'hefd,
12'heaa,
12'he5a,
12'he5b,
12'hea9,
12'hefe,
12'hf19,
12'hee7,
12'hea7,
12'he99,
12'hea5,
12'heca,
12'hf14,
12'hf68,
12'hf76,
12'hf27,
12'hece,
12'hebc,
12'hf00,
12'hf6a,
12'hfb6,
12'hfcb,
12'hfc2,
12'hfa7,
12'hf85,
12'hf70,
12'hf7f,
12'hfa9,
12'hfc3,
12'hfb6,
12'hf9b,
12'hfa4,
12'hfd9,
12'h01c,
12'h069,
12'h0b7,
12'h0e1,
12'h0e3,
12'h0bc,
12'h09a,
12'h0ab,
12'h0dd,
12'h114,
12'h135,
12'h13b,
12'h124,
12'h0fa,
12'h0dd,
12'h0e4,
12'h110,
12'h143,
12'h155,
12'h13e,
12'h108,
12'h0d4,
12'h0a1,
12'h06e,
12'h056,
12'h06a,
12'h0a3,
12'h0dd,
12'h0f4,
12'h0d5,
12'h0a7,
12'h095,
12'h0a4,
12'h0b6,
12'h0ab,
12'h08b,
12'h054,
12'h002,
12'hfaa,
12'hf74,
12'hf90,
12'hfe0,
12'hffe,
12'hfd2,
12'hf7e,
12'hf24,
12'hed6,
12'heb1,
12'heca,
12'heee,
12'hee4,
12'he91,
12'he38,
12'he1d,
12'he41,
12'he8f,
12'heda,
12'hf0c,
12'hf06,
12'heba,
12'he69,
12'he59,
12'he81,
12'hea2,
12'hea1,
12'hea3,
12'hed6,
12'hf14,
12'hf22,
12'hf27,
12'hf47,
12'hf6a,
12'hf4c,
12'hee0,
12'he85,
12'he69,
12'he83,
12'he8f,
12'he69,
12'he59,
12'he9b,
12'hf14,
12'hf70,
12'hf88,
12'hf6d,
12'hf35,
12'heee,
12'hec2,
12'hedd,
12'hf37,
12'hf90,
12'hf8f,
12'hf57,
12'hf5a,
12'hfb2,
12'h02a,
12'h06e,
12'h042,
12'hfc6,
12'hf44,
12'hf05,
12'hf31,
12'hfc3,
12'h07c,
12'h0ff,
12'h119,
12'h0d6,
12'h07e,
12'h073,
12'h0d8,
12'h170,
12'h1cf,
12'h1c3,
12'h165,
12'h0fb,
12'h0e1,
12'h14d,
12'h220,
12'h2fe,
12'h381,
12'h37e,
12'h317,
12'h2b0,
12'h296,
12'h2b5,
12'h2d1,
12'h2be,
12'h277,
12'h204,
12'h180,
12'h144,
12'h189,
12'h21b,
12'h27f,
12'h262,
12'h1fd,
12'h19d,
12'h15e,
12'h151,
12'h172,
12'h18e,
12'h160,
12'h0d6,
12'h037,
12'hfe8,
12'h01c,
12'h09d,
12'h0e7,
12'h0c3,
12'h041,
12'hfb1,
12'hf80,
12'hfc2,
12'h013,
12'h026,
12'hfdb,
12'hf40,
12'hea6,
12'he56,
12'he84,
12'hf10,
12'hf83,
12'hf87,
12'hf2e,
12'hec5,
12'he8b,
12'he95,
12'hee3,
12'hf36,
12'hf47,
12'hf10,
12'heb6,
12'he7e,
12'he85,
12'hea7,
12'heb9,
12'hec0,
12'heb2,
12'he8f,
12'he7a,
12'he94,
12'hede,
12'hf26,
12'hf4b,
12'hf3d,
12'heff,
12'hed8,
12'hf0c,
12'hf91,
12'hff9,
12'hff2,
12'hfa8,
12'hf50,
12'hf1a,
12'hf1f,
12'hf4d,
12'hf82,
12'hf9b,
12'hf8f,
12'hf6a,
12'hf4d,
12'hf65,
12'hfb8,
12'h029,
12'h08a,
12'h096,
12'h069,
12'h045,
12'h052,
12'h093,
12'h0eb,
12'h13e,
12'h170,
12'h161,
12'h122,
12'h0e6,
12'h0cc,
12'h0ea,
12'h112,
12'h129,
12'h131,
12'h12d,
12'h120,
12'h10e,
12'h0f8,
12'h0cd,
12'h08d,
12'h05c,
12'h05a,
12'h088,
12'h0c8,
12'h0ef,
12'h0ef,
12'h0df,
12'h0d2,
12'h0b4,
12'h08d,
12'h068,
12'h03c,
12'h005,
12'hfc9,
12'hf9c,
12'hf9a,
12'hfc6,
12'h000,
12'h028,
12'h018,
12'hfb8,
12'hf24,
12'hea7,
12'he80,
12'heb0,
12'hef1,
12'hf03,
12'hee1,
12'heb0,
12'he91,
12'he89,
12'he91,
12'hea8,
12'hebb,
12'hea8,
12'he6a,
12'he30,
12'he23,
12'he4d,
12'heb6,
12'hf2c,
12'hf65,
12'hf59,
12'hf2d,
12'hf02,
12'heed,
12'hef0,
12'hefc,
12'hf17,
12'hf2e,
12'hf05,
12'he8f,
12'he18,
12'hded,
12'he1d,
12'he8c,
12'hf00,
12'hf4f,
12'hf85,
12'hfab,
12'hfb9,
12'hfbd,
12'hfd7,
12'hfea,
12'hfad,
12'hf33,
12'heba,
12'he77,
12'he7e,
12'hebb,
12'hf3c,
12'hfe7,
12'h072,
12'h0b3,
12'h0a0,
12'h069,
12'h02f,
12'hfe9,
12'hfae,
12'hfa3,
12'hfd0,
12'hff9,
12'h011,
12'h053,
12'h0e6,
12'h1a4,
12'h22b,
12'h243,
12'h215,
12'h1ed,
12'h1bb,
12'h17d,
12'h170,
12'h1b5,
12'h219,
12'h252,
12'h25d,
12'h274,
12'h2ac,
12'h2d8,
12'h2df,
12'h2c3,
12'h2a3,
12'h270,
12'h23a,
12'h232,
12'h240,
12'h242,
12'h226,
12'h1f3,
12'h1b4,
12'h171,
12'h141,
12'h13f,
12'h16c,
12'h18f,
12'h16f,
12'h124,
12'h0e1,
12'h0a9,
12'h075,
12'h05c,
12'h060,
12'h05f,
12'h049,
12'h02f,
12'h023,
12'h023,
12'h007,
12'hfaf,
12'hf31,
12'hecf,
12'head,
12'heb9,
12'hed1,
12'hefc,
12'hf41,
12'hf92,
12'hfbb,
12'hf9f,
12'hf73,
12'hf56,
12'hf33,
12'heea,
12'he80,
12'he39,
12'he2b,
12'he46,
12'he72,
12'he9e,
12'hecd,
12'heea,
12'hed3,
12'he90,
12'he62,
12'he77,
12'hec3,
12'hf12,
12'hf4c,
12'hf60,
12'hf3c,
12'hefe,
12'hed0,
12'hed5,
12'hf1e,
12'hf88,
12'hfc5,
12'hfb5,
12'hf82,
12'hf72,
12'hf95,
12'hfc0,
12'hfd0,
12'hfb5,
12'hf88,
12'hf52,
12'hf1d,
12'hf2c,
12'hf84,
12'hff2,
12'h045,
12'h06c,
12'h083,
12'h08d,
12'h08d,
12'h092,
12'h0ce,
12'h133,
12'h16b,
12'h156,
12'h11c,
12'h0f7,
12'h0e8,
12'h0d7,
12'h0d3,
12'h0fc,
12'h141,
12'h16d,
12'h15f,
12'h127,
12'h0d5,
12'h08a,
12'h075,
12'h098,
12'h0cd,
12'h0ea,
12'h0e7,
12'h0d3,
12'h0b8,
12'h095,
12'h078,
12'h072,
12'h06a,
12'h040,
12'hffb,
12'hfc2,
12'hfb3,
12'hfc0,
12'hfd2,
12'hfe8,
12'hff9,
12'hfda,
12'hf91,
12'hf62,
12'hf6b,
12'hf77,
12'hf5f,
12'hf1f,
12'hed5,
12'he98,
12'he5b,
12'he32,
12'he2e,
12'he54,
12'he91,
12'heb5,
12'heaa,
12'he86,
12'he67,
12'he51,
12'he30,
12'he16,
12'he28,
12'he56,
12'he81,
12'hea1,
12'hebb,
12'heef,
12'hf3e,
12'hf7d,
12'hf9b,
12'hf7e,
12'hf34,
12'hed9,
12'he8c,
12'he6f,
12'he6a,
12'he7d,
12'hea2,
12'hed4,
12'hf30,
12'hfaa,
12'h00b,
12'h031,
12'h00c,
12'hfbe,
12'hf6f,
12'hf1f,
12'hee4,
12'hec5,
12'heb8,
12'hec0,
12'hee2,
12'hf35,
12'hfca,
12'h085,
12'h11e,
12'h139,
12'h0d5,
12'h055,
12'hff9,
12'hfdc,
12'hff2,
12'h018,
12'h041,
12'h04f,
12'h05a,
12'h099,
12'h135,
12'h20e,
12'h2b4,
12'h2d2,
12'h284,
12'h203,
12'h191,
12'h155,
12'h144,
12'h17e,
12'h1ed,
12'h248,
12'h25e,
12'h271,
12'h2be,
12'h31d,
12'h34c,
12'h326,
12'h2c9,
12'h246,
12'h1be,
12'h170,
12'h18a,
12'h1d9,
12'h20d,
12'h1f6,
12'h1a5,
12'h158,
12'h136,
12'h14b,
12'h171,
12'h190,
12'h174,
12'h110,
12'h08e,
12'h025,
12'h00c,
12'h036,
12'h072,
12'h079,
12'h038,
12'hfe3,
12'hfa0,
12'hf78,
12'hf7e,
12'hf98,
12'hf79,
12'hf04,
12'he7c,
12'he35,
12'he3f,
12'he92,
12'hf15,
12'hf8d,
12'hfba,
12'hf85,
12'hf2b,
12'hefb,
12'hef7,
12'heea,
12'heb3,
12'he73,
12'he4d,
12'he45,
12'he49,
12'he5f,
12'he98,
12'hed1,
12'heea,
12'hede,
12'hece,
12'hee5,
12'hf11,
12'hf3e,
12'hf62,
12'hf68,
12'hf44,
12'hf00,
12'hedc,
12'hf08,
12'hf6e,
12'hfc0,
12'hfe4,
12'hfe0,
12'hfc1,
12'hfb1,
12'hfc6,
12'hfe4,
12'hfeb,
12'hfe4,
12'hfd7,
12'hfb8,
12'hf8c,
12'hf9d,
12'h00d,
12'h08b,
12'h0bf,
12'h0b2,
12'h0ab,
12'h0ba,
12'h0b4,
12'h09f,
12'h0ae,
12'h0fc,
12'h167,
12'h198,
12'h180,
12'h151,
12'h11d,
12'h0ef,
12'h0cc,
12'h0d4,
12'h125,
12'h175,
12'h174,
12'h135,
12'h0ed,
12'h0be,
12'h09e,
12'h096,
12'h0be,
12'h0ef,
12'h0f3,
12'h0c8,
12'h093,
12'h07b,
12'h07e,
12'h080,
12'h07d,
12'h055,
12'h00a,
12'hfba,
12'hf7f,
12'hf81,
12'hfac,
12'hfe3,
12'h003,
12'hfe6,
12'hf9b,
12'hf4f,
12'hf17,
12'hefb,
12'hedc,
12'hebc,
12'he9a,
12'he67,
12'he37,
12'he18,
12'he2c,
12'he7d,
12'hed1,
12'hed8,
12'he9a,
12'he6f,
12'he71,
12'he71,
12'he4c,
12'he36,
12'he5e,
12'he9d,
12'hea9,
12'he8f,
12'heaa,
12'hf01,
12'hf4b,
12'hf5d,
12'hf3a,
12'hf02,
12'hecd,
12'he86,
12'he3f,
12'he19,
12'he23,
12'he4d,
12'he88,
12'hef7,
12'hf8f,
12'h00a,
12'h03f,
12'h023,
12'hfdc,
12'hf93,
12'hf53,
12'hf18,
12'hee2,
12'hec7,
12'hed9,
12'hf14,
12'hf5c,
12'hfae,
12'h016,
12'h089,
12'h0c3,
12'h0b6,
12'h08d,
12'h05f,
12'h033,
12'hffa,
12'hfcc,
12'hfd4,
12'h00b,
12'h04b,
12'h0a1,
12'h127,
12'h1b0,
12'h201,
12'h210,
12'h213,
12'h231,
12'h23e,
12'h202,
12'h1ae,
12'h1a2,
12'h1f1,
12'h251,
12'h284,
12'h2ac,
12'h2f7,
12'h33b,
12'h31d,
12'h2bf,
12'h269,
12'h22f,
12'h21b,
12'h212,
12'h1fd,
12'h1de,
12'h1a8,
12'h177,
12'h172,
12'h187,
12'h188,
12'h16e,
12'h152,
12'h14a,
12'h137,
12'h10e,
12'h0e4,
12'h0be,
12'h094,
12'h058,
12'h01f,
12'hff9,
12'hff9,
12'h00f,
12'h00f,
12'hfe5,
12'hf9d,
12'hf47,
12'heea,
12'hea4,
12'he93,
12'heb3,
12'hed6,
12'heeb,
12'hf00,
12'hf20,
12'hf38,
12'hf35,
12'hf2f,
12'hf2e,
12'hf22,
12'hee1,
12'he72,
12'he2b,
12'he45,
12'he98,
12'hed1,
12'hecf,
12'hec0,
12'hec6,
12'heca,
12'heab,
12'he96,
12'hebf,
12'hf02,
12'hf3d,
12'hf5c,
12'hf58,
12'hf30,
12'hef9,
12'hedd,
12'heeb,
12'hf20,
12'hf56,
12'hf6c,
12'hf63,
12'hf67,
12'hf95,
12'hfd6,
12'hff9,
12'hffc,
12'hff9,
12'hfe2,
12'hfa8,
12'hf6e,
12'hf8f,
12'hffc,
12'h066,
12'h0a4,
12'h0b0,
12'h0b5,
12'h0b4,
12'h094,
12'h07d,
12'h0ae,
12'h11b,
12'h189,
12'h19c,
12'h153,
12'h104,
12'h0d3,
12'h0c7,
12'h0e2,
12'h122,
12'h166,
12'h170,
12'h132,
12'h0d5,
12'h08f,
12'h090,
12'h0c5,
12'h0ed,
12'h0ee,
12'h0c8,
12'h0a3,
12'h096,
12'h099,
12'h0b2,
12'h0c1,
12'h0af,
12'h07f,
12'h044,
12'h01c,
12'h013,
12'h016,
12'h013,
12'h007,
12'hfe3,
12'hfaf,
12'hf77,
12'hf4b,
12'hf43,
12'hf48,
12'hf34,
12'hf02,
12'hed3,
12'heb9,
12'hea3,
12'he8d,
12'he89,
12'hea8,
12'hedd,
12'hef1,
12'hed9,
12'hebe,
12'heaf,
12'heb4,
12'he9e,
12'he5e,
12'he34,
12'he3f,
12'he77,
12'hebf,
12'hf01,
12'hf3f,
12'hf77,
12'hf85,
12'hf4e,
12'hef9,
12'hebd,
12'he9f,
12'he7f,
12'he5e,
12'he53,
12'he77,
12'heaf,
12'hed0,
12'heff,
12'hf59,
12'hfb7,
12'hfe7,
12'hfdc,
12'hfae,
12'hf6d,
12'hf1a,
12'hed0,
12'hebc,
12'hed6,
12'hefc,
12'hf21,
12'hf4f,
12'hf95,
12'hff4,
12'h063,
12'h0a7,
12'h09d,
12'h061,
12'h00b,
12'hfb1,
12'hf7d,
12'hf83,
12'hfbf,
12'h00a,
12'h03e,
12'h077,
12'h0d6,
12'h155,
12'h1bc,
12'h1f3,
12'h204,
12'h1e8,
12'h1b6,
12'h16a,
12'h124,
12'h134,
12'h1b3,
12'h257,
12'h2c0,
12'h2ea,
12'h301,
12'h31f,
12'h325,
12'h2f1,
12'h291,
12'h216,
12'h197,
12'h148,
12'h149,
12'h184,
12'h1ce,
12'h1ff,
12'h20a,
12'h1fc,
12'h1da,
12'h1a4,
12'h170,
12'h15a,
12'h148,
12'h117,
12'h0d0,
12'h07b,
12'h042,
12'h036,
12'h048,
12'h05d,
12'h061,
12'h05b,
12'h03e,
12'h014,
12'hff9,
12'hfe9,
12'hfbf,
12'hf62,
12'hef5,
12'heb5,
12'heaa,
12'hebf,
12'hef1,
12'hf46,
12'hf8f,
12'hf89,
12'hf56,
12'hf41,
12'hf54,
12'hf4e,
12'hef3,
12'he78,
12'he41,
12'he4d,
12'he6d,
12'he9a,
12'hed6,
12'hf19,
12'hf38,
12'hf1e,
12'hef7,
12'hf02,
12'hf2d,
12'hf4a,
12'hf5c,
12'hf60,
12'hf42,
12'hf01,
12'hed5,
12'hef3,
12'hf60,
12'hfc7,
12'hfed,
12'hfd9,
12'hfa5,
12'hf7b,
12'hf79,
12'hfa9,
12'hfd8,
12'hff2,
12'hff9,
12'hfd8,
12'hf98,
12'hf72,
12'hf9d,
12'h014,
12'h08d,
12'h0bf,
12'h0b9,
12'h097,
12'h06a,
12'h04d,
12'h071,
12'h0ce,
12'h13b,
12'h162,
12'h12d,
12'h0e2,
12'h0c9,
12'h0db,
12'h0e8,
12'h0ff,
12'h126,
12'h139,
12'h10a,
12'h0ae,
12'h058,
12'h044,
12'h064,
12'h080,
12'h086,
12'h085,
12'h09b,
12'h0bf,
12'h0da,
12'h0d0,
12'h0b0,
12'h08d,
12'h060,
12'h029,
12'hfef,
12'hfce,
12'hfc7,
12'hfce,
12'hfd4,
12'hfd5,
12'hfda,
12'hfcf,
12'hfa9,
12'hf76,
12'hf44,
12'hf18,
12'hee7,
12'heb2,
12'he9b,
12'he95,
12'he8a,
12'he6e,
12'he6f,
12'heb3,
12'hef4,
12'hef5,
12'hec6,
12'he9e,
12'he94,
12'he94,
12'he7a,
12'he52,
12'he4a,
12'he67,
12'he8d,
12'hea2,
12'hec2,
12'hf14,
12'hf6b,
12'hf9f,
12'hf9e,
12'hf72,
12'hf3a,
12'hee8,
12'he84,
12'he43,
12'he3f,
12'he5b,
12'he6e,
12'he89,
12'hee6,
12'hf7f,
12'hffc,
12'h015,
12'hfd9,
12'hf8f,
12'hf49,
12'hf04,
12'hed5,
12'hecd,
12'hef0,
12'hf14,
12'hf31,
12'hf75,
12'hff6,
12'h08a,
12'h0da,
12'h0c4,
12'h07e,
12'h028,
12'hfda,
12'hfb4,
12'hfd0,
12'h019,
12'h054,
12'h055,
12'h03d,
12'h066,
12'h0e9,
12'h192,
12'h20d,
12'h22c,
12'h20b,
12'h1bc,
12'h15f,
12'h127,
12'h140,
12'h1bb,
12'h252,
12'h29f,
12'h296,
12'h288,
12'h2bc,
12'h314,
12'h343,
12'h328,
12'h2b3,
12'h20e,
12'h184,
12'h154,
12'h186,
12'h1e6,
12'h227,
12'h228,
12'h1fb,
12'h1c6,
12'h1a6,
12'h1a1,
12'h1aa,
12'h19b,
12'h160,
12'h0ee,
12'h079,
12'h033,
12'h03b,
12'h075,
12'h097,
12'h080,
12'h044,
12'h001,
12'hfd3,
12'hfdd,
12'h00b,
12'h00b,
12'hf9e,
12'heee,
12'he64,
12'he47,
12'he7b,
12'hecf,
12'hf31,
12'hf73,
12'hf68,
12'hf19,
12'hede,
12'hef3,
12'hf2a,
12'hf2c,
12'hecb,
12'he50,
12'he1f,
12'he32,
12'he5c,
12'he89,
12'heba,
12'hee7,
12'hed7,
12'he9f,
12'he92,
12'hed3,
12'hf2a,
12'hf4b,
12'hf45,
12'hf2b,
12'hef0,
12'heae,
12'hea8,
12'hf07,
12'hf8c,
12'hfcb,
12'hfb1,
12'hf80,
12'hf70,
12'hf8a,
12'hfc1,
12'hfeb,
12'hfe9,
12'hfcb,
12'hf94,
12'hf4c,
12'hf33,
12'hf88,
12'h022,
12'h098,
12'h0b5,
12'h09a,
12'h083,
12'h086,
12'h086,
12'h092,
12'h0cd,
12'h11b,
12'h151,
12'h148,
12'h11f,
12'h10e,
12'h10d,
12'h108,
12'h0f1,
12'h0f5,
12'h124,
12'h13e,
12'h128,
12'h0f6,
12'h0ca,
12'h0b4,
12'h0a2,
12'h08c,
12'h095,
12'h0ba,
12'h0da,
12'h0d4,
12'h0b9,
12'h0ac,
12'h0ac,
12'h0ad,
12'h09a,
12'h071,
12'h033,
12'hffc,
12'hfdc,
12'hfcb,
12'hfe5,
12'h025,
12'h046,
12'h028,
12'hfd8,
12'hf7f,
12'hf34,
12'hef3,
12'hedb,
12'hee0,
12'hee1,
12'hebd,
12'he82,
12'he6e,
12'he9b,
12'hee5,
12'hf07,
12'hee8,
12'heb0,
12'he83,
12'he66,
12'he5d,
12'he6a,
12'he94,
12'hebd,
12'hec3,
12'heb1,
12'hea4,
12'hec8,
12'hf10,
12'hf5c,
12'hf9e,
12'hfaf,
12'hf7b,
12'hf19,
12'heae,
12'he63,
12'he59,
12'he7f,
12'hea1,
12'hea0,
12'he8f,
12'heaa,
12'hf12,
12'hf98,
12'hfe5,
12'hfdb,
12'hf90,
12'hf0a,
12'he8d,
12'he64,
12'hea4,
12'hf14,
12'hf55,
12'hf6c,
12'hf97,
12'h001,
12'h086,
12'h0d5,
12'h0d1,
12'h07f,
12'hff9,
12'hf7a,
12'hf4a,
12'hf8a,
12'h003,
12'h064,
12'h099,
12'h0c1,
12'h0ff,
12'h155,
12'h1a8,
12'h1d8,
12'h1e2,
12'h1a8,
12'h12b,
12'h0b4,
12'h0b1,
12'h154,
12'h243,
12'h2f3,
12'h323,
12'h308,
12'h2e8,
12'h2df,
12'h2e8,
12'h2f9,
12'h2e4,
12'h28a,
12'h1fd,
12'h174,
12'h126,
12'h13a,
12'h19a,
12'h1fc,
12'h224,
12'h1f6,
12'h1a2,
12'h171,
12'h181,
12'h1a6,
12'h1a3,
12'h15d,
12'h0e4,
12'h05c,
12'hfed,
12'hfd4,
12'h007,
12'h045,
12'h06e,
12'h072,
12'h054,
12'h02a,
12'h00f,
12'hffc,
12'hfbb,
12'hf54,
12'hee1,
12'he84,
12'he61,
12'he8a,
12'hefc,
12'hf7d,
12'hfc2,
12'hfa0,
12'hf4e,
12'hf1b,
12'hf12,
12'hefb,
12'hebe,
12'he83,
12'he6b,
12'he69,
12'he71,
12'he8d,
12'hec6,
12'hef7,
12'hef4,
12'hebf,
12'he96,
12'heb8,
12'hf0c,
12'hf58,
12'hf83,
12'hf84,
12'hf4c,
12'heed,
12'hea5,
12'heb6,
12'hf16,
12'hf82,
12'hfbe,
12'hfbc,
12'hfa8,
12'hfa9,
12'hfd4,
12'h001,
12'hfff,
12'hfd1,
12'hf89,
12'hf3c,
12'hf13,
12'hf47,
12'hfe1,
12'h08d,
12'h0ef,
12'h0fc,
12'h0d6,
12'h092,
12'h056,
12'h05d,
12'h0af,
12'h107,
12'h126,
12'h103,
12'h0c9,
12'h0c7,
12'h100,
12'h140,
12'h15d,
12'h15f,
12'h158,
12'h132,
12'h0ed,
12'h0a2,
12'h084,
12'h09a,
12'h0a7,
12'h09c,
12'h07d,
12'h072,
12'h09c,
12'h0c9,
12'h0d6,
12'h0ab,
12'h075,
12'h060,
12'h04e,
12'h028,
12'hff5,
12'hfd4,
12'hfcd,
12'hfb6,
12'hf8c,
12'hf89,
12'hfb4,
12'hfe0,
12'hfe7,
12'hfce,
12'hf93,
12'hf33,
12'hecc,
12'he97,
12'he9c,
12'he88,
12'he52,
12'he29,
12'he32,
12'he6f,
12'heb5,
12'hedb,
12'hee8,
12'hef0,
12'hee3,
12'heaa,
12'he6e,
12'he73,
12'heaf,
12'hee5,
12'hee6,
12'hec8,
12'heba,
12'heda,
12'hf1a,
12'hf5f,
12'hf7f,
12'hf6b,
12'hf27,
12'hebf,
12'he61,
12'he2a,
12'he33,
12'he63,
12'head,
12'hf0b,
12'hf60,
12'hfa7,
12'hfd9,
12'hfff,
12'h013,
12'h00e,
12'hfdd,
12'hf6f,
12'hef1,
12'heaa,
12'hebe,
12'heff,
12'hf3b,
12'hf7d,
12'hfdd,
12'h03f,
12'h070,
12'h060,
12'h03c,
12'h023,
12'h009,
12'hff0,
12'hff1,
12'h004,
12'h009,
12'h00d,
12'h045,
12'h0cb,
12'h182,
12'h21f,
12'h25d,
12'h245,
12'h20f,
12'h1d7,
12'h18f,
12'h15e,
12'h199,
12'h218,
12'h272,
12'h281,
12'h29e,
12'h2ea,
12'h325,
12'h322,
12'h2df,
12'h28f,
12'h23a,
12'h1e1,
12'h1ac,
12'h1b8,
12'h1e9,
12'h202,
12'h1f3,
12'h1cc,
12'h196,
12'h15d,
12'h153,
12'h17d,
12'h1ae,
12'h1a9,
12'h152,
12'h0dc,
12'h07a,
12'h053,
12'h06c,
12'h091,
12'h094,
12'h062,
12'h00f,
12'hfc7,
12'hfa8,
12'hfb0,
12'hfb1,
12'hf81,
12'hf20,
12'heb5,
12'he76,
12'he74,
12'head,
12'hf16,
12'hf8d,
12'hfc8,
12'hf9f,
12'hf41,
12'hf02,
12'hf00,
12'hf01,
12'hed9,
12'he96,
12'he76,
12'he71,
12'he69,
12'he6c,
12'he96,
12'heec,
12'hf1d,
12'hefc,
12'heb1,
12'he92,
12'hec1,
12'hf0a,
12'hf3c,
12'hf53,
12'hf41,
12'hf06,
12'hec9,
12'hec8,
12'hf16,
12'hf78,
12'hfb5,
12'hfbb,
12'hfa3,
12'hf89,
12'hf90,
12'hfae,
12'hfd0,
12'hfdd,
12'hfc9,
12'hf8f,
12'hf53,
12'hf5b,
12'hfae,
12'h018,
12'h057,
12'h06d,
12'h077,
12'h07d,
12'h077,
12'h087,
12'h0ce,
12'h131,
12'h176,
12'h16d,
12'h12c,
12'h0e8,
12'h0c2,
12'h0c4,
12'h0da,
12'h0ff,
12'h137,
12'h158,
12'h147,
12'h108,
12'h0c2,
12'h0a0,
12'h09e,
12'h0a5,
12'h0b8,
12'h0d0,
12'h0e0,
12'h0e8,
12'h0dc,
12'h0b6,
12'h082,
12'h058,
12'h03d,
12'h022,
12'hff8,
12'hfde,
12'hfe1,
12'hfe5,
12'hfe2,
12'hfea,
12'hff7,
12'hfd0,
12'hf77,
12'hf31,
12'hf22,
12'hf21,
12'hf07,
12'hee7,
12'hedc,
12'hec6,
12'he8f,
12'he68,
12'he75,
12'heaa,
12'hed7,
12'hed5,
12'heb4,
12'he8f,
12'he81,
12'he74,
12'he54,
12'he4b,
12'he6f,
12'heaa,
12'hed1,
12'hed9,
12'hee1,
12'hf09,
12'hf4b,
12'hf87,
12'hf90,
12'hf53,
12'hefc,
12'hea8,
12'he67,
12'he54,
12'he6d,
12'he8f,
12'he9d,
12'hec5,
12'hf27,
12'hfa1,
12'hff8,
12'hff4,
12'hfb6,
12'hf61,
12'hf10,
12'hece,
12'he9e,
12'he96,
12'heb2,
12'heec,
12'hf28,
12'hf7c,
12'hff3,
12'h071,
12'h0c5,
12'h0b8,
12'h068,
12'h004,
12'hfc0,
12'hfb1,
12'hfcf,
12'h006,
12'h039,
12'h057,
12'h07f,
12'h0d5,
12'h156,
12'h1c2,
12'h1e1,
12'h1c2,
12'h195,
12'h174,
12'h168,
12'h168,
12'h192,
12'h1fb,
12'h264,
12'h298,
12'h2a1,
12'h2cd,
12'h323,
12'h355,
12'h330,
12'h2d2,
12'h270,
12'h21d,
12'h1e3,
12'h1cd,
12'h1df,
12'h1fc,
12'h205,
12'h1fb,
12'h1eb,
12'h1da,
12'h1c6,
12'h1ac,
12'h193,
12'h169,
12'h119,
12'h0b4,
12'h05b,
12'h032,
12'h049,
12'h078,
12'h086,
12'h07e,
12'h07c,
12'h074,
12'h05d,
12'h039,
12'hffe,
12'hf8f,
12'hef2,
12'he76,
12'he69,
12'heae,
12'hefc,
12'hf43,
12'hf8c,
12'hfb5,
12'hf99,
12'hf54,
12'hf2c,
12'hf30,
12'hf1b,
12'hebb,
12'he3d,
12'he04,
12'he25,
12'he5c,
12'he8d,
12'heb6,
12'hed9,
12'hede,
12'heba,
12'hea2,
12'hec9,
12'hf1d,
12'hf58,
12'hf5c,
12'hf3f,
12'hf0f,
12'hed0,
12'he94,
12'hea1,
12'hf02,
12'hf6d,
12'hf9c,
12'hf8e,
12'hf79,
12'hf6e,
12'hf80,
12'hf94,
12'hf9b,
12'hfa6,
12'hfa8,
12'hf95,
12'hf6e,
12'hf72,
12'hfcf,
12'h05e,
12'h0cc,
12'h0e2,
12'h0bc,
12'h088,
12'h04f,
12'h030,
12'h04a,
12'h0ab,
12'h128,
12'h16d,
12'h15b,
12'h11f,
12'h0ef,
12'h0cf,
12'h0ce,
12'h0f5,
12'h13b,
12'h16f,
12'h157,
12'h0fc,
12'h09a,
12'h079,
12'h087,
12'h08e,
12'h095,
12'h0a8,
12'h0b4,
12'h09d,
12'h07f,
12'h07f,
12'h093,
12'h0a3,
12'h08b,
12'h051,
12'h000,
12'hfbb,
12'hfa9,
12'hfc0,
12'hfe8,
12'h008,
12'h018,
12'hff1,
12'hf9b,
12'hf5b,
12'hf4c,
12'hf53,
12'hf35,
12'heeb,
12'he98,
12'he60,
12'he52,
12'he5b,
12'he78,
12'hea5,
12'hec8,
12'hec5,
12'he9b,
12'he8b,
12'heb1,
12'hedf,
12'hed3,
12'he9a,
12'he78,
12'he89,
12'hebb,
12'hedb,
12'heed,
12'hf18,
12'hf49,
12'hf68,
12'hf5b,
12'hf33,
12'hf12,
12'hef0,
12'heae,
12'he64,
12'he3e,
12'he36,
12'he44,
12'he84,
12'hf10,
12'hfa8,
12'hff9,
12'hff3,
12'hfb9,
12'hf85,
12'hf54,
12'hf22,
12'hef7,
12'hec7,
12'hea5,
12'heac,
12'heec,
12'hf64,
12'hffc,
12'h084,
12'h0c9,
12'h0ba,
12'h07d,
12'h040,
12'h011,
12'hff6,
12'hfe0,
12'hfce,
12'hfbc,
12'hfbc,
12'hffc,
12'h099,
12'h169,
12'h1f7,
12'h214,
12'h1d8,
12'h1a7,
12'h1b5,
12'h1d1,
12'h1dd,
12'h1dc,
12'h1ef,
12'h218,
12'h22e,
12'h245,
12'h2a1,
12'h338,
12'h38c,
12'h351,
12'h2c1,
12'h22b,
12'h1c0,
12'h1ae,
12'h1ec,
12'h22e,
12'h233,
12'h1e9,
12'h199,
12'h18a,
12'h196,
12'h1a2,
12'h1ae,
12'h1b0,
12'h187,
12'h121,
12'h0c3,
12'h0a5,
12'h0b8,
12'h0c6,
12'h0ac,
12'h06f,
12'h02a,
12'h010,
12'h024,
12'h050,
12'h06e,
12'h040,
12'hfb4,
12'heed,
12'he50,
12'he34,
12'he89,
12'hef6,
12'hf4b,
12'hf8d,
12'hf9f,
12'hf6e,
12'hf2e,
12'hf20,
12'hf40,
12'hf3e,
12'heea,
12'he5e,
12'he0c,
12'he22,
12'he73,
12'hec0,
12'hef9,
12'hf19,
12'hf00,
12'hebc,
12'he7b,
12'he8b,
12'hef2,
12'hf54,
12'hf77,
12'hf6d,
12'hf4d,
12'hf0b,
12'hec2,
12'heb1,
12'heee,
12'hf41,
12'hf6e,
12'hf7b,
12'hf81,
12'hf91,
12'hfbc,
12'hfe5,
12'hfde,
12'hfb8,
12'hfa5,
12'hf98,
12'hf72,
12'hf61,
12'hf9c,
12'h013,
12'h074,
12'h08e,
12'h082,
12'h07a,
12'h06d,
12'h03b,
12'h018,
12'h053,
12'h0dd,
12'h14c,
12'h162,
12'h143,
12'h11e,
12'h0f7,
12'h0d0,
12'h0bf,
12'h0e9,
12'h125,
12'h128,
12'h0e6,
12'h087,
12'h05f,
12'h07b,
12'h0a8,
12'h0c4,
12'h0c8,
12'h0b0,
12'h07d,
12'h05a,
12'h062,
12'h087,
12'h0a9,
12'h0af,
12'h085,
12'h034,
12'hfed,
12'hfd0,
12'hfdd,
12'h000,
12'h024,
12'h028,
12'hff4,
12'hf93,
12'hf40,
12'hf27,
12'hf3a,
12'hf3d,
12'hf09,
12'heba,
12'he78,
12'he60,
12'he64,
12'he78,
12'heba,
12'hf0f,
12'hf31,
12'hf0a,
12'hecd,
12'heb6,
12'hec0,
12'heaa,
12'he72,
12'he59,
12'he70,
12'he97,
12'heb0,
12'hece,
12'hf1d,
12'hf81,
12'hfb2,
12'hf8c,
12'hf31,
12'hef5,
12'hed5,
12'he9f,
12'he58,
12'he38,
12'he48,
12'he69,
12'hea1,
12'hf1b,
12'hfbe,
12'h018,
12'h006,
12'hfba,
12'hf72,
12'hf4b,
12'hf2f,
12'hf19,
12'hefd,
12'hee2,
12'hee3,
12'hf0a,
12'hf64,
12'hfde,
12'h05e,
12'h0b0,
12'h0a6,
12'h073,
12'h044,
12'h01b,
12'hffd,
12'hfdb,
12'hfc1,
12'hfc4,
12'hfd9,
12'h00c,
12'h08d,
12'h14d,
12'h1fc,
12'h251,
12'h248,
12'h221,
12'h1f9,
12'h1c9,
12'h18a,
12'h161,
12'h18e,
12'h201,
12'h25a,
12'h274,
12'h29d,
12'h2e9,
12'h327,
12'h31f,
12'h2cf,
12'h267,
12'h1fd,
12'h1bf,
12'h1c8,
12'h1fc,
12'h230,
12'h237,
12'h20c,
12'h1d4,
12'h1a0,
12'h171,
12'h153,
12'h159,
12'h173,
12'h160,
12'h12a,
12'h0f9,
12'h0c3,
12'h096,
12'h081,
12'h069,
12'h056,
12'h03a,
12'h010,
12'hff8,
12'hff5,
12'hff5,
12'hfc9,
12'hf65,
12'hef3,
12'heaf,
12'heaf,
12'hed8,
12'hf12,
12'hf67,
12'hfab,
12'hf9c,
12'hf48,
12'hefe,
12'hef2,
12'hefb,
12'hed4,
12'he7b,
12'he34,
12'he29,
12'he5b,
12'he98,
12'hec5,
12'hef6,
12'hf18,
12'hf01,
12'heb7,
12'he8b,
12'he9d,
12'hed2,
12'hf00,
12'hf1b,
12'hf28,
12'hf16,
12'heef,
12'hed5,
12'hefb,
12'hf49,
12'hf81,
12'hf90,
12'hf78,
12'hf64,
12'hf74,
12'hf9a,
12'hfaf,
12'hfb9,
12'hfbf,
12'hfae,
12'hf76,
12'hf46,
12'hf74,
12'hfe7,
12'h055,
12'h089,
12'h09c,
12'h0af,
12'h0a5,
12'h07f,
12'h063,
12'h090,
12'h105,
12'h169,
12'h17a,
12'h143,
12'h104,
12'h0df,
12'h0ca,
12'h0c8,
12'h0f2,
12'h12d,
12'h12e,
12'h0ed,
12'h0a0,
12'h079,
12'h085,
12'h09e,
12'h0ad,
12'h0b1,
12'h0ae,
12'h0b0,
12'h0bf,
12'h0cf,
12'h0dd,
12'h0d8,
12'h0b1,
12'h071,
12'h01e,
12'hfe4,
12'hfd5,
12'hfd9,
12'hfe9,
12'hffc,
12'h00b,
12'h002,
12'hfcf,
12'hf8b,
12'hf52,
12'hf2d,
12'hf11,
12'hef1,
12'hee1,
12'hee1,
12'hed8,
12'heac,
12'he82,
12'he8e,
12'hec6,
12'heed,
12'hed3,
12'he94,
12'he60,
12'he63,
12'he71,
12'he67,
12'he6a,
12'he8d,
12'heb3,
12'hebb,
12'hec3,
12'heef,
12'hf49,
12'hf98,
12'hfa7,
12'hf77,
12'hf2b,
12'hee6,
12'hea8,
12'he77,
12'he6a,
12'he84,
12'he9a,
12'hea1,
12'hed3,
12'hf38,
12'hfb6,
12'h002,
12'hffa,
12'hfbe,
12'hf5e,
12'hef5,
12'heb9,
12'hece,
12'hf10,
12'hf4c,
12'hf6e,
12'hf8f,
12'hfe9,
12'h06f,
12'h0e4,
12'h10a,
12'h0dd,
12'h087,
12'h017,
12'hfb1,
12'hf8b,
12'hfa6,
12'hfdc,
12'h017,
12'h050,
12'h0a8,
12'h12f,
12'h1bc,
12'h21e,
12'h238,
12'h219,
12'h1d2,
12'h179,
12'h133,
12'h125,
12'h168,
12'h1ef,
12'h268,
12'h297,
12'h2a9,
12'h2e0,
12'h33b,
12'h370,
12'h351,
12'h2e8,
12'h25c,
12'h1e0,
12'h191,
12'h17b,
12'h1a5,
12'h1e6,
12'h1f7,
12'h1d4,
12'h1a7,
12'h195,
12'h1a2,
12'h1b8,
12'h1b5,
12'h193,
12'h155,
12'h0e6,
12'h069,
12'h019,
12'h011,
12'h02c,
12'h03e,
12'h03e,
12'h033,
12'h02d,
12'h034,
12'h045,
12'h030,
12'hfd0,
12'hf20,
12'he7c,
12'he52,
12'he8d,
12'heeb,
12'hf41,
12'hf77,
12'hf66,
12'hf13,
12'hed2,
12'hedd,
12'hf13,
12'hf25,
12'hef8,
12'he90,
12'he33,
12'he32,
12'he73,
12'hece,
12'hf0f,
12'hf14,
12'hecb,
12'he6b,
12'he53,
12'hea0,
12'hf20,
12'hf67,
12'hf72,
12'hf53,
12'hf07,
12'hea6,
12'he6d,
12'heb1,
12'hf33,
12'hf7b,
12'hf6b,
12'hf4b,
12'hf52,
12'hf8c,
12'hfdf,
12'hfff,
12'hfeb,
12'hfc1,
12'hf8e,
12'hf4b,
12'hf22,
12'hf67,
12'hff5,
12'h078,
12'h0b0,
12'h0a3,
12'h091,
12'h08a,
12'h082,
12'h088,
12'h0c2,
12'h113,
12'h140,
12'h135,
12'h110,
12'h106,
12'h11b,
12'h131,
12'h12c,
12'h11a,
12'h10e,
12'h0ed,
12'h0c0,
12'h0a5,
12'h0a3,
12'h0b7,
12'h0c4,
12'h0b4,
12'h09e,
12'h0a0,
12'h0ac,
12'h0a9,
12'h092,
12'h082,
12'h083,
12'h082,
12'h07b,
12'h059,
12'h022,
12'hff2,
12'hfcc,
12'hfb4,
12'hfa5,
12'hf9f,
12'hfa7,
12'hfb9,
12'hfb3,
12'hf8c,
12'hf5b,
12'hf2c,
12'hf06,
12'hedd,
12'heab,
12'he64,
12'he21,
12'he10,
12'he45,
12'hea0,
12'hee2,
12'heee,
12'hec1,
12'he8f,
12'he88,
12'he90,
12'he8a,
12'he89,
12'he9a,
12'heb0,
12'hec2,
12'hec9,
12'heef,
12'hf3d,
12'hf84,
12'hfa2,
12'hf73,
12'hf22,
12'hee0,
12'he99,
12'he60,
12'he55,
12'he79,
12'he98,
12'he9e,
12'hebb,
12'hf17,
12'hf96,
12'hfd6,
12'hfc2,
12'hf91,
12'hf55,
12'hf13,
12'hef8,
12'hf14,
12'hf39,
12'hf51,
12'hf57,
12'hf59,
12'hf90,
12'h012,
12'h088,
12'h09f,
12'h075,
12'h03b,
12'hffe,
12'hfcf,
12'hfc1,
12'hfcc,
12'hfe3,
12'h000,
12'h02e,
12'h084,
12'h115,
12'h1bc,
12'h224,
12'h233,
12'h211,
12'h1d3,
12'h193,
12'h15a,
12'h149,
12'h183,
12'h1e5,
12'h259,
12'h2b3,
12'h2e5,
12'h31f,
12'h349,
12'h339,
12'h2f8,
12'h28b,
12'h211,
12'h1b5,
12'h189,
12'h19a,
12'h1d7,
12'h20d,
12'h222,
12'h20c,
12'h1dd,
12'h1b6,
12'h18a,
12'h15c,
12'h13c,
12'h122,
12'h0fc,
12'h0c4,
12'h088,
12'h061,
12'h05a,
12'h065,
12'h05d,
12'h043,
12'h023,
12'hffb,
12'hfee,
12'hfed,
12'hfc7,
12'hf69,
12'hef3,
12'heab,
12'he9c,
12'heaa,
12'hec3,
12'hef7,
12'hf3b,
12'hf4f,
12'hf2d,
12'hf11,
12'hf20,
12'hf2d,
12'hef1,
12'he84,
12'he38,
12'he3c,
12'he6e,
12'he9e,
12'hebf,
12'hee1,
12'hefd,
12'hef0,
12'hed1,
12'hedb,
12'hf07,
12'hf26,
12'hf1f,
12'hf11,
12'hf0d,
12'hf06,
12'heed,
12'hee0,
12'hf17,
12'hf7f,
12'hfc0,
12'hfb2,
12'hf97,
12'hfa0,
12'hfcc,
12'hff9,
12'h000,
12'hffd,
12'hffc,
12'hfec,
12'hfab,
12'hf63,
12'hf75,
12'hfde,
12'h05b,
12'h0a3,
12'h0bb,
12'h0c1,
12'h0b9,
12'h0a9,
12'h0aa,
12'h0e6,
12'h144,
12'h17d,
12'h16f,
12'h138,
12'h110,
12'h108,
12'h105,
12'h0fe,
12'h110,
12'h131,
12'h140,
12'h118,
12'h0b7,
12'h074,
12'h080,
12'h0a9,
12'h0b8,
12'h0b8,
12'h0bd,
12'h0c1,
12'h0b3,
12'h0a5,
12'h0b5,
12'h0c6,
12'h0b4,
12'h067,
12'hffc,
12'hfbb,
12'hfb3,
12'hfc1,
12'hfca,
12'hfd3,
12'hfd7,
12'hfc9,
12'hfa5,
12'hf7a,
12'hf5e,
12'hf45,
12'hf11,
12'hed3,
12'heb2,
12'hea4,
12'he97,
12'he81,
12'he72,
12'he8a,
12'hec0,
12'hee7,
12'heda,
12'hea8,
12'he87,
12'he86,
12'he74,
12'he4b,
12'he39,
12'he5a,
12'he93,
12'heb1,
12'heb9,
12'hedb,
12'hf22,
12'hf66,
12'hf8c,
12'hf83,
12'hf45,
12'hefd,
12'heb6,
12'he5e,
12'he25,
12'he23,
12'he48,
12'he99,
12'hf17,
12'hfad,
12'h01a,
12'h029,
12'hfea,
12'hf8f,
12'hf45,
12'hf16,
12'hefb,
12'hef2,
12'hef8,
12'hf15,
12'hf45,
12'hf90,
12'h00f,
12'h09c,
12'h0e3,
12'h0da,
12'h098,
12'h03b,
12'hff4,
12'hfbe,
12'hfa2,
12'hfbf,
12'hff3,
12'h015,
12'h04a,
12'h0bf,
12'h169,
12'h1ff,
12'h242,
12'h23f,
12'h22a,
12'h219,
12'h1eb,
12'h19f,
12'h174,
12'h197,
12'h1ed,
12'h237,
12'h26b,
12'h2ba,
12'h31d,
12'h35a,
12'h349,
12'h2f3,
12'h289,
12'h21b,
12'h1cb,
12'h1b7,
12'h1c9,
12'h1ee,
12'h1f7,
12'h1dd,
12'h1c4,
12'h1ab,
12'h18c,
12'h16a,
12'h15a,
12'h15b,
12'h14c,
12'h122,
12'h0e0,
12'h09d,
12'h069,
12'h041,
12'h02a,
12'h028,
12'h028,
12'h01d,
12'h00a,
12'hff7,
12'hfd9,
12'hf8d,
12'hf14,
12'heb9,
12'heac,
12'hec5,
12'hecf,
12'hed3,
12'hf0b,
12'hf55,
12'hf5b,
12'hf2c,
12'hf0a,
12'hf10,
12'hf0a,
12'hebb,
12'he4f,
12'he30,
12'he61,
12'he9e,
12'hec4,
12'hed3,
12'hee3,
12'hee0,
12'heb9,
12'he84,
12'he81,
12'heca,
12'hf20,
12'hf40,
12'hf33,
12'hf17,
12'heed,
12'hec7,
12'hec8,
12'hf07,
12'hf58,
12'hf7d,
12'hf89,
12'hf94,
12'hfb1,
12'hfe6,
12'h001,
12'hfed,
12'hfcc,
12'hfb1,
12'hf82,
12'hf3f,
12'hf1b,
12'hf53,
12'hfdf,
12'h050,
12'h077,
12'h080,
12'h094,
12'h0a2,
12'h093,
12'h095,
12'h0d9,
12'h142,
12'h181,
12'h174,
12'h13f,
12'h117,
12'h104,
12'h0f4,
12'h0fc,
12'h11b,
12'h139,
12'h127,
12'h0d5,
12'h089,
12'h083,
12'h0ab,
12'h0d4,
12'h0d8,
12'h0bd,
12'h09e,
12'h083,
12'h087,
12'h0a5,
12'h0ca,
12'h0d9,
12'h0a9,
12'h040,
12'hfe4,
12'hfbc,
12'hfc3,
12'hfd2,
12'hfcd,
12'hfc7,
12'hfc3,
12'hfb9,
12'hf9d,
12'hf85,
12'hf7a,
12'hf57,
12'hf09,
12'heb3,
12'he87,
12'he8a,
12'he9a,
12'he97,
12'he91,
12'hea9,
12'hecf,
12'hed3,
12'heb3,
12'he99,
12'he99,
12'he8e,
12'he52,
12'he1b,
12'he2a,
12'he7d,
12'hec9,
12'hedb,
12'hee9,
12'hf27,
12'hf6f,
12'hf8d,
12'hf78,
12'hf50,
12'hf2c,
12'hefc,
12'heb3,
12'he64,
12'he3a,
12'he3e,
12'he59,
12'he9d,
12'hf35,
12'hfdb,
12'h01d,
12'hfef,
12'hf8f,
12'hf54,
12'hf39,
12'hf27,
12'hf20,
12'hf1e,
12'hf17,
12'hf12,
12'hf28,
12'hf89,
12'h034,
12'h0d3,
12'h107,
12'h0c9,
12'h06a,
12'h016,
12'hfcf,
12'hf9c,
12'hf96,
12'hfc3,
12'hff4,
12'h012,
12'h04d,
12'h0dc,
12'h19e,
12'h241,
12'h28e,
12'h27c,
12'h22a,
12'h1c5,
12'h157,
12'h100,
12'h108,
12'h180,
12'h218,
12'h279,
12'h2a8,
12'h2db,
12'h31e,
12'h339,
12'h316,
12'h2d1,
12'h275,
12'h20d,
12'h1bf,
12'h1a4,
12'h1ba,
12'h1e1,
12'h1e7,
12'h1d4,
12'h1af,
12'h171,
12'h12b,
12'h111,
12'h144,
12'h17d,
12'h173,
12'h127,
12'h0b7,
12'h051,
12'h01a,
12'h016,
12'h03b,
12'h052,
12'h041,
12'h012,
12'hfe4,
12'hfd9,
12'hfd4,
12'hfaf,
12'hf6c,
12'hf1c,
12'hed0,
12'he8f,
12'he6f,
12'hea0,
12'hf1a,
12'hf77,
12'hf67,
12'hf21,
12'hf06,
12'hf16,
12'hf0c,
12'hec8,
12'he84,
12'he78,
12'he82,
12'he80,
12'he85,
12'hea5,
12'hed9,
12'hef3,
12'hece,
12'hea2,
12'heb2,
12'heef,
12'hf22,
12'hf3a,
12'hf49,
12'hf4b,
12'hf1e,
12'hee1,
12'hef3,
12'hf50,
12'hfac,
12'hfd2,
12'hfcf,
12'hfc0,
12'hfc0,
12'hfd7,
12'hfe5,
12'hfda,
12'hfc9,
12'hfb0,
12'hf76,
12'hf31,
12'hf31,
12'hfa2,
12'h02e,
12'h074,
12'h086,
12'h09a,
12'h0be,
12'h0ce,
12'h0b9,
12'h0c0,
12'h10a,
12'h16b,
12'h18e,
12'h154,
12'h0fd,
12'h0d1,
12'h0cb,
12'h0cf,
12'h0ed,
12'h12d,
12'h160,
12'h150,
12'h108,
12'h0c6,
12'h0a5,
12'h09b,
12'h089,
12'h076,
12'h07b,
12'h09a,
12'h0c1,
12'h0df,
12'h0f1,
12'h0e4,
12'h0bb,
12'h07a,
12'h02a,
12'hff4,
12'hfe2,
12'hfde,
12'hfd0,
12'hfc7,
12'hfdc,
12'hffc,
12'h000,
12'hfe1,
12'hfab,
12'hf6d,
12'hf34,
12'hf06,
12'hef1,
12'heee,
12'hee5,
12'hec0,
12'he76,
12'he3f,
12'he5e,
12'hea0,
12'heba,
12'he9f,
12'he83,
12'he88,
12'he8e,
12'he74,
12'he5c,
12'he7e,
12'hec5,
12'hee3,
12'hed4,
12'hecb,
12'hef7,
12'hf40,
12'hf6c,
12'hf6e,
12'hf54,
12'hf3d,
12'hf0f,
12'heb9,
12'he69,
12'he3c,
12'he3d,
12'he5b,
12'heb1,
12'hf4b,
12'hfd1,
12'h00a,
12'hfff,
12'hfd1,
12'hfaf,
12'hf8e,
12'hf58,
12'hf22,
12'hef8,
12'hee7,
12'hf01,
12'hf48,
12'hfbe,
12'h047,
12'h0bb,
12'h0e1,
12'h0b0,
12'h06d,
12'h02d,
12'hfea,
12'hfac,
12'hf91,
12'hfb4,
12'hff6,
12'h04a,
12'h0bc,
12'h145,
12'h1bf,
12'h1fb,
12'h1ff,
12'h1f0,
12'h1eb,
12'h1dd,
12'h1a1,
12'h155,
12'h149,
12'h194,
12'h20d,
12'h272,
12'h2af,
12'h2e2,
12'h307,
12'h2ff,
12'h2ca,
12'h291,
12'h263,
12'h22c,
12'h1fe,
12'h1e6,
12'h1d2,
12'h1ba,
12'h1a6,
12'h1b0,
12'h1bb,
12'h19c,
12'h15e,
12'h12a,
12'h133,
12'h150,
12'h142,
12'h108,
12'h0b2,
12'h050,
12'hffa,
12'hfd7,
12'hff1,
12'h01f,
12'h043,
12'h04e,
12'h031,
12'hfeb,
12'hf88,
12'hf1a,
12'heac,
12'he62,
12'he55,
12'he68,
12'he87,
12'hec5,
12'hf2e,
12'hf83,
12'hf8b,
12'hf59,
12'hf1a,
12'hef1,
12'hecb,
12'he83,
12'he40,
12'he46,
12'he7e,
12'heac,
12'hebc,
12'hec4,
12'hed9,
12'hee6,
12'hec6,
12'hea0,
12'heb9,
12'hf00,
12'hf34,
12'hf3f,
12'hf3f,
12'hf38,
12'hf1e,
12'hef5,
12'heee,
12'hf21,
12'hf5e,
12'hf8c,
12'hfb4,
12'hfdb,
12'hff9,
12'hffb,
12'hfdf,
12'hfc5,
12'hfb5,
12'hfa7,
12'hf77,
12'hf33,
12'hf2e,
12'hf92,
12'h024,
12'h08e,
12'h0bb,
12'h0cc,
12'h0bf,
12'h088,
12'h05f,
12'h085,
12'h0f7,
12'h16f,
12'h1a0,
12'h17a,
12'h128,
12'h0eb,
12'h0da,
12'h0ef,
12'h11d,
12'h147,
12'h143,
12'h10b,
12'h0c2,
12'h09f,
12'h0b7,
12'h0e3,
12'h0f5,
12'h0e7,
12'h0d9,
12'h0d9,
12'h0e9,
12'h0f6,
12'h0f6,
12'h0e1,
12'h0b6,
12'h080,
12'h047,
12'h01f,
12'h012,
12'h00f,
12'h003,
12'hff2,
12'hfec,
12'hff3,
12'hfe4,
12'hfb7,
12'hf80,
12'hf54,
12'hf29,
12'heed,
12'heb7,
12'hea0,
12'he97,
12'he84,
12'he69,
12'he6d,
12'heaa,
12'hee3,
12'hee0,
12'heb8,
12'he98,
12'he93,
12'he88,
12'he5c,
12'he2d,
12'he25,
12'he46,
12'he72,
12'heb1,
12'hf06,
12'hf4d,
12'hf77,
12'hf89,
12'hf80,
12'hf62,
12'hf36,
12'hf02,
12'hec1,
12'he7f,
12'he61,
12'he7a,
12'heaa,
12'hee2,
12'hf30,
12'hf8c,
12'hfd3,
12'hfeb,
12'hfe0,
12'hfb2,
12'hf52,
12'hedb,
12'he8e,
12'he9b,
12'hef0,
12'hf47,
12'hf7c,
12'hfac,
12'h002,
12'h06a,
12'h0aa,
12'h0b6,
12'h097,
12'h04c,
12'hfdb,
12'hf7c,
12'hf70,
12'hfb2,
12'h005,
12'h037,
12'h060,
12'h0ad,
12'h11e,
12'h196,
12'h1f1,
12'h225,
12'h223,
12'h1ce,
12'h147,
12'h0e4,
12'h0f7,
12'h17e,
12'h21e,
12'h289,
12'h2bc,
12'h2eb,
12'h323,
12'h342,
12'h337,
12'h305,
12'h2aa,
12'h22e,
12'h1b3,
12'h164,
12'h162,
12'h197,
12'h1db,
12'h216,
12'h219,
12'h1f2,
12'h1cf,
12'h1be,
12'h1bb,
12'h19d,
12'h159,
12'h103,
12'h09e,
12'h04a,
12'h01b,
12'h023,
12'h046,
12'h051,
12'h039,
12'h009,
12'hff1,
12'hff6,
12'hff8,
12'hfd0,
12'hf6a,
12'heed,
12'he86,
12'he50,
12'he5b,
12'heb0,
12'hf25,
12'hf65,
12'hf50,
12'hf19,
12'hf08,
12'hf24,
12'hf35,
12'hf0a,
12'hea5,
12'he50,
12'he18,
12'he08,
12'he35,
12'he92,
12'hef8,
12'hf21,
12'hef6,
12'heb9,
12'hec2,
12'hf08,
12'hf3c,
12'hf4b,
12'hf51,
12'hf49,
12'hf0e,
12'heb4,
12'he97,
12'heec,
12'hf7c,
12'hfd3,
12'hfd3,
12'hfad,
12'hf8e,
12'hf94,
12'hfbb,
12'hfe5,
12'hffa,
12'hff1,
12'hfba,
12'hf6d,
12'hf56,
12'hf96,
12'h00c,
12'h07d,
12'h0c6,
12'h0d3,
12'h0ae,
12'h06f,
12'h04a,
12'h07c,
12'h0e9,
12'h14b,
12'h159,
12'h11f,
12'h0e7,
12'h0d8,
12'h0f3,
12'h10e,
12'h115,
12'h117,
12'h115,
12'h10b,
12'h0f5,
12'h0d9,
12'h0ca,
12'h0c3,
12'h0a7,
12'h068,
12'h036,
12'h048,
12'h092,
12'h0c9,
12'h0db,
12'h0d8,
12'h0d6,
12'h0d9,
12'h0af,
12'h053,
12'hff5,
12'hfaa,
12'hf7b,
12'hf74,
12'hf9e,
12'hfe1,
12'h003,
12'hff3,
12'hfca,
12'hf98,
12'hf51,
12'hef2,
12'heab,
12'he9d,
12'he9c,
12'he93,
12'he87,
12'he8a,
12'heb3,
12'hed9,
12'hede,
12'hec0,
12'he9a,
12'he97,
12'heaa,
12'heba,
12'hebf,
12'hed0,
12'heec,
12'heef,
12'heda,
12'hebf,
12'hec7,
12'hefb,
12'hf33,
12'hf54,
12'hf5e,
12'hf64,
12'hf5d,
12'hf1e,
12'heb9,
12'he69,
12'he4d,
12'he52,
12'he75,
12'hed5,
12'hf57,
12'hfc3,
12'hff5,
12'hff5,
12'hfdc,
12'hfac,
12'hf6f,
12'hf36,
12'hf05,
12'hee4,
12'hedb,
12'hefc,
12'hf5d,
12'hff1,
12'h087,
12'h0d7,
12'h0bf,
12'h073,
12'h02b,
12'hff8,
12'hfd4,
12'hfb5,
12'hfb6,
12'hfd7,
12'hfec,
12'h005,
12'h067,
12'h115,
12'h1bc,
12'h209,
12'h1f5,
12'h1c3,
12'h1be,
12'h1d1,
12'h1c9,
12'h1c5,
12'h1eb,
12'h225,
12'h243,
12'h245,
12'h270,
12'h2c6,
12'h309,
12'h301,
12'h2ae,
12'h256,
12'h20d,
12'h1e0,
12'h1e7,
12'h209,
12'h21e,
12'h1f7,
12'h1aa,
12'h176,
12'h16d,
12'h173,
12'h165,
12'h164,
12'h16d,
12'h150,
12'h112,
12'h0cc,
12'h0a2,
12'h0a0,
12'h094,
12'h064,
12'h028,
12'h005,
12'h005,
12'h017,
12'h032,
12'h03c,
12'hfef,
12'hf38,
12'he6e,
12'he1d,
12'he5c,
12'heb5,
12'hef8,
12'hf40,
12'hf87,
12'hf94,
12'hf54,
12'hf23,
12'hf30,
12'hf38,
12'heed,
12'he51,
12'hddb,
12'hde5,
12'he3d,
12'hea1,
12'hee9,
12'hf06,
12'hef5,
12'heae,
12'he62,
12'he54,
12'he8d,
12'hede,
12'hf0a,
12'hf1c,
12'hf2a,
12'hf16,
12'hee1,
12'hec0,
12'hee0,
12'hf26,
12'hf4f,
12'hf50,
12'hf56,
12'hf73,
12'hfad,
12'hfeb,
12'h00e,
12'h012,
12'hfef,
12'hfb1,
12'hf5e,
12'hf20,
12'hf3c,
12'hfb5,
12'h041,
12'h096,
12'h0a9,
12'h0a5,
12'h0b0,
12'h0b5,
12'h0af,
12'h0c1,
12'h105,
12'h157,
12'h166,
12'h13b,
12'h116,
12'h109,
12'h10e,
12'h111,
12'h11c,
12'h12a,
12'h123,
12'h0ec,
12'h094,
12'h068,
12'h083,
12'h0be,
12'h0ed,
12'h0ff,
12'h0f1,
12'h0d0,
12'h099,
12'h064,
12'h063,
12'h08a,
12'h0aa,
12'h098,
12'h04e,
12'h008,
12'hfec,
12'hff1,
12'hff9,
12'hfeb,
12'hfd0,
12'hfb0,
12'hf8a,
12'hf63,
12'hf5b,
12'hf73,
12'hf7d,
12'hf50,
12'hefc,
12'hebb,
12'he91,
12'he78,
12'he71,
12'he8a,
12'hec2,
12'hef5,
12'hf02,
12'hef5,
12'hef3,
12'hef4,
12'heca,
12'he81,
12'he4e,
12'he57,
12'he9c,
12'hedc,
12'hf03,
12'hf33,
12'hf6d,
12'hf8b,
12'hf71,
12'hf3d,
12'hf21,
12'hf1d,
12'hef9,
12'he9c,
12'he41,
12'he2a,
12'he5e,
12'heb9,
12'hf35,
12'hfc6,
12'h02a,
12'h027,
12'hfcd,
12'hf74,
12'hf5d,
12'hf6f,
12'hf71,
12'hf48,
12'hf03,
12'hec9,
12'heb8,
12'heea,
12'hf69,
12'h01e,
12'h0c1,
12'h0ed,
12'h0a7,
12'h03f,
12'hff1,
12'hfd6,
12'hfe5,
12'h00c,
12'h025,
12'h00c,
12'hfde,
12'h001,
12'h0b1,
12'h1ab,
12'h272,
12'h2b3,
12'h27d,
12'h20c,
12'h19a,
12'h14f,
12'h152,
12'h1ab,
12'h220,
12'h254,
12'h236,
12'h227,
12'h26a,
12'h2da,
12'h32a,
12'h334,
12'h2e0,
12'h242,
12'h1a5,
12'h16f,
12'h1ba,
12'h22a,
12'h252,
12'h21a,
12'h1d0,
12'h196,
12'h164,
12'h156,
12'h17d,
12'h1b0,
12'h199,
12'h12b,
12'h0aa,
12'h05d,
12'h064,
12'h097,
12'h0bf,
12'h0b7,
12'h06e,
12'h002,
12'hfb0,
12'hfa4,
12'hfcd,
12'hfe5,
12'hfac,
12'hf3a,
12'hecb,
12'he87,
12'he7b,
12'hea1,
12'hee6,
12'hf2d,
12'hf5b,
12'hf47,
12'heff,
12'hed4,
12'heeb,
12'hf0a,
12'hef1,
12'heaa,
12'he69,
12'he34,
12'he12,
12'he18,
12'he55,
12'head,
12'hee0,
12'hed2,
12'heaf,
12'heb9,
12'hee2,
12'hf10,
12'hf2f,
12'hf37,
12'hf1d,
12'heec,
12'hec1,
12'hec0,
12'hf09,
12'hf67,
12'hf9a,
12'hf95,
12'hf82,
12'hf85,
12'hf92,
12'hf8e,
12'hf84,
12'hf91,
12'hfa1,
12'hf93,
12'hf74,
12'hf7c,
12'hfc6,
12'h012,
12'h037,
12'h04e,
12'h073,
12'h0b3,
12'h0d1,
12'h0b5,
12'h0b1,
12'h0e5,
12'h123,
12'h135,
12'h120,
12'h106,
12'h0ec,
12'h0c0,
12'h09b,
12'h0b3,
12'h111,
12'h167,
12'h167,
12'h115,
12'h0ac,
12'h060,
12'h042,
12'h053,
12'h092,
12'h0d4,
12'h0ed,
12'h0d9,
12'h0b1,
12'h094,
12'h089,
12'h093,
12'h093,
12'h074,
12'h041,
12'h006,
12'hfd6,
12'hfba,
12'hfca,
12'h004,
12'h02b,
12'h011,
12'hfbb,
12'hf60,
12'hf35,
12'hf2f,
12'hf30,
12'hf28,
12'hf1c,
12'hef2,
12'hea5,
12'he52,
12'he45,
12'he9c,
12'hefb,
12'hf15,
12'hee7,
12'hea4,
12'he82,
12'he73,
12'he63,
12'he69,
12'hea3,
12'hee5,
12'hefe,
12'hee1,
12'hed1,
12'hf07,
12'hf4b,
12'hf66,
12'hf4b,
12'hf1b,
12'hef3,
12'hec5,
12'he8b,
12'he66,
12'he6a,
12'he81,
12'heaa,
12'hef8,
12'hf67,
12'hfdc,
12'h022,
12'h015,
12'hfdd,
12'hfb2,
12'hf96,
12'hf6b,
12'hf1e,
12'hed7,
12'hebf,
12'hecc,
12'hef5,
12'hf5e,
12'h006,
12'h0af,
12'h0fe,
12'h0da,
12'h085,
12'h022,
12'hfce,
12'hfa8,
12'hfbd,
12'h000,
12'h032,
12'h02c,
12'h025,
12'h080,
12'h13d,
12'h1fd,
12'h25b,
12'h24c,
12'h204,
12'h1b7,
12'h173,
12'h142,
12'h157,
12'h1c0,
12'h23a,
12'h25f,
12'h24b,
12'h26e,
12'h2c8,
12'h31c,
12'h32f,
12'h2f3,
12'h28e,
12'h222,
12'h1d7,
12'h1c1,
12'h1d5,
12'h1e6,
12'h1d1,
12'h1a5,
12'h178,
12'h146,
12'h12a,
12'h143,
12'h187,
12'h1b8,
12'h186,
12'h101,
12'h06d,
12'h017,
12'h01e,
12'h04c,
12'h06b,
12'h066,
12'h03c,
12'h000,
12'hfd3,
12'hfd2,
12'hfdc,
12'hfaf,
12'hf3c,
12'heb4,
12'he58,
12'he43,
12'he6d,
12'hed1,
12'hf5a,
12'hfbd,
12'hfaf,
12'hf4a,
12'hef4,
12'hee1,
12'hef1,
12'hee5,
12'heac,
12'he81,
12'he7d,
12'he6e,
12'he4e,
12'he50,
12'he96,
12'hed8,
12'hec3,
12'he7d,
12'he6e,
12'heb7,
12'hf20,
12'hf67,
12'hf7c,
12'hf65,
12'hf12,
12'heac,
12'he88,
12'hece,
12'hf3b,
12'hf7b,
12'hf82,
12'hf81,
12'hf8c,
12'hfa3,
12'hfb7,
12'hfb8,
12'hfba,
12'hfb3,
12'hf8a,
12'hf55,
12'hf50,
12'hfa2,
12'h020,
12'h071,
12'h07b,
12'h071,
12'h081,
12'h087,
12'h074,
12'h082,
12'h0d3,
12'h13a,
12'h168,
12'h145,
12'h104,
12'h0df,
12'h0d5,
12'h0d4,
12'h0e8,
12'h10c,
12'h12e,
12'h13c,
12'h118,
12'h0d1,
12'h0a6,
12'h0a5,
12'h0ae,
12'h0b9,
12'h0c1,
12'h0bf,
12'h0bd,
12'h0b4,
12'h09f,
12'h090,
12'h092,
12'h098,
12'h084,
12'h061,
12'h033,
12'hffc,
12'hfcf,
12'hfbb,
12'hfba,
12'hfcf,
12'hfe3,
12'hfcc,
12'hf9a,
12'hf6e,
12'hf50,
12'hf41,
12'hf34,
12'hf18,
12'hef6,
12'hebf,
12'he82,
12'he6f,
12'hea0,
12'heef,
12'hf14,
12'hefe,
12'hec5,
12'hea0,
12'he96,
12'he85,
12'he63,
12'he6d,
12'hea5,
12'hed5,
12'hee4,
12'heec,
12'hf10,
12'hf3c,
12'hf50,
12'hf34,
12'hf03,
12'hee2,
12'heca,
12'heaf,
12'he93,
12'he85,
12'he8f,
12'he9c,
12'heb2,
12'hf02,
12'hf8d,
12'hffc,
12'h010,
12'hfd5,
12'hf7c,
12'hf33,
12'hf0a,
12'hf06,
12'hf10,
12'hf19,
12'hf10,
12'hf01,
12'hf25,
12'hfa4,
12'h052,
12'h0d8,
12'h0eb,
12'h095,
12'h022,
12'hfb6,
12'hf75,
12'hf87,
12'hfdd,
12'h03c,
12'h058,
12'h041,
12'h059,
12'h0d8,
12'h199,
12'h231,
12'h26c,
12'h24e,
12'h1e2,
12'h15c,
12'h0ed,
12'h0dd,
12'h13e,
12'h1d9,
12'h268,
12'h2a1,
12'h2a4,
12'h2b7,
12'h2e7,
12'h315,
12'h31b,
12'h2f0,
12'h291,
12'h205,
12'h190,
12'h180,
12'h1bb,
12'h1fe,
12'h218,
12'h1f9,
12'h1b0,
12'h15b,
12'h13a,
12'h167,
12'h1b3,
12'h1cf,
12'h18f,
12'h10c,
12'h075,
12'h027,
12'h046,
12'h091,
12'h0c0,
12'h0a7,
12'h051,
12'hfea,
12'hfaf,
12'hfae,
12'hfbe,
12'hf9e,
12'hf39,
12'hed2,
12'he95,
12'he7a,
12'he9b,
12'hf01,
12'hf7b,
12'hfaf,
12'hf6c,
12'hefb,
12'heb8,
12'heb9,
12'hec3,
12'hea2,
12'he71,
12'he59,
12'he53,
12'he46,
12'he3d,
12'he5e,
12'heab,
12'hedb,
12'hece,
12'heb8,
12'hec4,
12'hee0,
12'heeb,
12'hef8,
12'hf14,
12'hf16,
12'hee4,
12'heaa,
12'hebc,
12'hf21,
12'hf85,
12'hfa8,
12'hfa0,
12'hf8f,
12'hf86,
12'hf8f,
12'hf91,
12'hf90,
12'hfaa,
12'hfb8,
12'hf8d,
12'hf50,
12'hf5c,
12'hfc9,
12'h047,
12'h08b,
12'h094,
12'h097,
12'h09b,
12'h093,
12'h097,
12'h0cb,
12'h12b,
12'h179,
12'h170,
12'h132,
12'h0fe,
12'h0f2,
12'h103,
12'h107,
12'h10b,
12'h127,
12'h14e,
12'h150,
12'h11c,
12'h0e4,
12'h0c4,
12'h0b6,
12'h0ac,
12'h0a9,
12'h0be,
12'h0e0,
12'h0fb,
12'h0fb,
12'h0e3,
12'h0d0,
12'h0c9,
12'h0b2,
12'h08e,
12'h062,
12'h03d,
12'h01c,
12'hff1,
12'hfd8,
12'hff2,
12'h020,
12'h015,
12'hfd6,
12'hf95,
12'hf65,
12'hf3e,
12'hf1e,
12'hf14,
12'hf10,
12'hef2,
12'heb1,
12'he72,
12'he6a,
12'hea2,
12'hed6,
12'hed8,
12'heb6,
12'hea3,
12'hea2,
12'he9b,
12'he8d,
12'he8c,
12'heb2,
12'hedf,
12'hee9,
12'heda,
12'hee7,
12'hf16,
12'hf3b,
12'hf4b,
12'hf3f,
12'hf13,
12'hedf,
12'hea5,
12'he6e,
12'he66,
12'he7b,
12'he78,
12'he61,
12'he79,
12'hee1,
12'hf76,
12'hfe3,
12'hff1,
12'hfb6,
12'hf5a,
12'hefb,
12'hebf,
12'hec0,
12'hef6,
12'hf25,
12'hf2b,
12'hf2d,
12'hf5c,
12'hfd6,
12'h063,
12'h0b7,
12'h0b2,
12'h06c,
12'h00a,
12'hfac,
12'hf77,
12'hf7f,
12'hfc5,
12'h01c,
12'h05b,
12'h08b,
12'h0db,
12'h15a,
12'h1e1,
12'h23b,
12'h255,
12'h235,
12'h1eb,
12'h184,
12'h13d,
12'h15d,
12'h1e4,
12'h28d,
12'h2ea,
12'h2de,
12'h2bd,
12'h2bf,
12'h2df,
12'h2ea,
12'h2d3,
12'h2a1,
12'h251,
12'h207,
12'h1d6,
12'h1cf,
12'h1ec,
12'h20c,
12'h20d,
12'h1dc,
12'h19b,
12'h162,
12'h150,
12'h166,
12'h185,
12'h190,
12'h161,
12'h0eb,
12'h06a,
12'h020,
12'h018,
12'h045,
12'h076,
12'h080,
12'h05b,
12'h01d,
12'hfec,
12'hfba,
12'hf71,
12'hf17,
12'hed3,
12'hebe,
12'hebb,
12'hec2,
12'hee7,
12'hf39,
12'hf82,
12'hf7a,
12'hf39,
12'hefd,
12'hed9,
12'heb0,
12'he65,
12'he26,
12'he30,
12'he72,
12'heaa,
12'hebf,
12'hec8,
12'hec8,
12'he9d,
12'he5b,
12'he49,
12'he8d,
12'hef1,
12'hf2b,
12'hf29,
12'hf16,
12'hf05,
12'hed4,
12'he9d,
12'heaf,
12'hf14,
12'hf72,
12'hf8d,
12'hf7e,
12'hf87,
12'hfbd,
12'hff5,
12'h009,
12'hfed,
12'hfc0,
12'hf83,
12'hf2f,
12'heeb,
12'hefa,
12'hf8a,
12'h041,
12'h0ae,
12'h0ae,
12'h087,
12'h079,
12'h077,
12'h08f,
12'h0da,
12'h141,
12'h186,
12'h176,
12'h129,
12'h0ee,
12'h0ee,
12'h107,
12'h10a,
12'h0f4,
12'h0e5,
12'h0e1,
12'h0d3,
12'h0b7,
12'h0b7,
12'h0d3,
12'h0ca,
12'h0a5,
12'h083,
12'h08d,
12'h0bb,
12'h0d6,
12'h0d7,
12'h0c8,
12'h0c4,
12'h0b9,
12'h08a,
12'h057,
12'h038,
12'h02e,
12'h01b,
12'hfe3,
12'hf9f,
12'hf84,
12'hf95,
12'hfa3,
12'hfaa,
12'hfbb,
12'hfb2,
12'hf6d,
12'hf07,
12'hebf,
12'heb9,
12'hec3,
12'hea9,
12'he70,
12'he4f,
12'he6c,
12'he96,
12'head,
12'hec4,
12'hee9,
12'hef8,
12'hec9,
12'he6f,
12'he2f,
12'he46,
12'he98,
12'hedf,
12'hf08,
12'hf1a,
12'hf1f,
12'hf15,
12'hf0d,
12'hf0d,
12'hf09,
12'hefb,
12'hecf,
12'he82,
12'he37,
12'he28,
12'he61,
12'hecc,
12'hf50,
12'hfb9,
12'hfef,
12'hfe6,
12'hfa2,
12'hf70,
12'hf78,
12'hf8b,
12'hf71,
12'hf1a,
12'hebb,
12'he9c,
12'hec2,
12'hef9,
12'hf59,
12'h008,
12'h0af,
12'h0d5,
12'h08e,
12'h042,
12'h033,
12'h050,
12'h053,
12'h032,
12'hffc,
12'hfd2,
12'hfcd,
12'h027,
12'h105,
12'h20f,
12'h2bd,
12'h2bc,
12'h24e,
12'h1eb,
12'h1c4,
12'h1ba,
12'h1c0,
12'h1e9,
12'h226,
12'h252,
12'h260,
12'h280,
12'h2e7,
12'h35e,
12'h382,
12'h337,
12'h29b,
12'h203,
12'h1ba,
12'h1d1,
12'h21f,
12'h25a,
12'h246,
12'h1f1,
12'h19d,
12'h170,
12'h162,
12'h174,
12'h18a,
12'h188,
12'h14f,
12'h0e7,
12'h095,
12'h077,
12'h089,
12'h0a2,
12'h096,
12'h055,
12'hff0,
12'hf9b,
12'hf8a,
12'hfbd,
12'hfef,
12'hfd3,
12'hf5a,
12'hec0,
12'he61,
12'he57,
12'he7a,
12'heba,
12'hf1a,
12'hf6d,
12'hf74,
12'hf22,
12'hed0,
12'hed5,
12'hefa,
12'hef9,
12'hea7,
12'he3d,
12'he15,
12'he17,
12'he29,
12'he53,
12'he99,
12'hed4,
12'hede,
12'heb3,
12'he89,
12'he9e,
12'hee5,
12'hf28,
12'hf4b,
12'hf5a,
12'hf52,
12'hf25,
12'hee1,
12'heca,
12'hefb,
12'hf46,
12'hf7a,
12'hf8f,
12'hfa1,
12'hfb1,
12'hfbb,
12'hfbb,
12'hfb5,
12'hfc0,
12'hfc6,
12'hfb2,
12'hfa3,
12'hfbe,
12'h001,
12'h037,
12'h04e,
12'h078,
12'h0d5,
12'h129,
12'h121,
12'h0da,
12'h0bf,
12'h108,
12'h173,
12'h1b0,
12'h1ae,
12'h18a,
12'h14b,
12'h0f3,
12'h0be,
12'h0da,
12'h139,
12'h18f,
12'h19d,
12'h165,
12'h118,
12'h0d0,
12'h0a9,
12'h0c6,
12'h101,
12'h128,
12'h112,
12'h0d3,
12'h0a3,
12'h09e,
12'h0c5,
12'h0f5,
12'h0f9,
12'h0bd,
12'h05a,
12'h006,
12'hfe1,
12'hfe9,
12'h003,
12'h01a,
12'h017,
12'hfdc,
12'hf8e,
12'hf58,
12'hf4c,
12'hf59,
12'hf4c,
12'hf0f,
12'hec4,
12'he8f,
12'he69,
12'he5b,
12'he7a,
12'hec4,
12'hef7,
12'hedf,
12'he84,
12'he32,
12'he20,
12'he3a,
12'he4e,
12'he5a,
12'he71,
12'he79,
12'he7a,
12'he84,
12'hebf,
12'hf28,
12'hf76,
12'hf71,
12'hf26,
12'hece,
12'he91,
12'he70,
12'he5b,
12'he58,
12'he61,
12'he56,
12'he4a,
12'he77,
12'hefa,
12'hf99,
12'hff4,
12'hfdd,
12'hf78,
12'hf18,
12'hed9,
12'hec4,
12'hed7,
12'heff,
12'hf1b,
12'hf23,
12'hf31,
12'hf79,
12'h01a,
12'h0bb,
12'h0fc,
12'h0da,
12'h081,
12'h00c,
12'hfae,
12'hf87,
12'hf8c,
12'hfb1,
12'hfe1,
12'h00d,
12'h051,
12'h0cb,
12'h171,
12'h20a,
12'h256,
12'h24b,
12'h207,
12'h1c2,
12'h181,
12'h156,
12'h174,
12'h1e2,
12'h26f,
12'h2b5,
12'h2be,
12'h2d8,
12'h2fb,
12'h31a,
12'h317,
12'h2e0,
12'h296,
12'h243,
12'h205,
12'h1e1,
12'h1db,
12'h1e9,
12'h1e7,
12'h1c3,
12'h180,
12'h146,
12'h126,
12'h133,
12'h162,
12'h185,
12'h189,
12'h155,
12'h0ec,
12'h07f,
12'h03f,
12'h035,
12'h032,
12'h021,
12'h00a,
12'hff0,
12'hfe1,
12'hfec,
12'hfe7,
12'hf9b,
12'hf1c,
12'heb4,
12'he8e,
12'he8b,
12'he9f,
12'hedb,
12'hf41,
12'hf7b,
12'hf5b,
12'hf10,
12'hedb,
12'hedb,
12'hed2,
12'he95,
12'he55,
12'he50,
12'he70,
12'he8f,
12'hea1,
12'heac,
12'heab,
12'he9a,
12'he81,
12'he7b,
12'heb3,
12'hefd,
12'hf32,
12'hf44,
12'hf42,
12'hf28,
12'hef6,
12'hec1,
12'hec8,
12'hf15,
12'hf52,
12'hf5e,
12'hf62,
12'hf80,
12'hfb7,
12'hfde,
12'hfd8,
12'hfbd,
12'hfa4,
12'hf7f,
12'hf3d,
12'hf0a,
12'hf2f,
12'hfa3,
12'h01e,
12'h07c,
12'h0a4,
12'h0b7,
12'h0b6,
12'h083,
12'h061,
12'h075,
12'h0d1,
12'h14c,
12'h189,
12'h172,
12'h13f,
12'h118,
12'h104,
12'h104,
12'h120,
12'h153,
12'h16c,
12'h13f,
12'h0e5,
12'h0aa,
12'h0a4,
12'h0b2,
12'h0c3,
12'h0d9,
12'h0e5,
12'h0dc,
12'h0bf,
12'h0a0,
12'h099,
12'h0aa,
12'h0b6,
12'h0a5,
12'h073,
12'h034,
12'h00b,
12'hfec,
12'hfc7,
12'hfb3,
12'hfc5,
12'hfe1,
12'hfdb,
12'hfbe,
12'hf99,
12'hf6d,
12'hf2b,
12'hede,
12'heab,
12'hea1,
12'he98,
12'he7a,
12'he5a,
12'he5b,
12'he93,
12'heca,
12'hed5,
12'hec0,
12'hea7,
12'he91,
12'he60,
12'he27,
12'he1c,
12'he4c,
12'he93,
12'hec3,
12'heda,
12'hf00,
12'hf24,
12'hf1d,
12'hef4,
12'hec2,
12'heb4,
12'heb8,
12'he9a,
12'he5a,
12'he24,
12'he21,
12'he57,
12'hec2,
12'hf49,
12'hfc5,
12'h005,
12'hff2,
12'hfa6,
12'hf6b,
12'hf5d,
12'hf69,
12'hf59,
12'hf1d,
12'hed6,
12'heac,
12'hecb,
12'hf28,
12'hfc3,
12'h072,
12'h0da,
12'h0c6,
12'h068,
12'h01d,
12'h016,
12'h03a,
12'h055,
12'h058,
12'h050,
12'h025,
12'h00a,
12'h067,
12'h143,
12'h23a,
12'h2b4,
12'h295,
12'h22e,
12'h1de,
12'h1b6,
12'h19c,
12'h1a5,
12'h1e8,
12'h246,
12'h264,
12'h24b,
12'h26d,
12'h2dd,
12'h346,
12'h35a,
12'h30e,
12'h280,
12'h1df,
12'h18f,
12'h1b0,
12'h20c,
12'h25b,
12'h252,
12'h1ff,
12'h1ad,
12'h177,
12'h166,
12'h18a,
12'h1ba,
12'h1c4,
12'h179,
12'h0f1,
12'h084,
12'h064,
12'h083,
12'h0a8,
12'h0a6,
12'h062,
12'hff3,
12'hf9f,
12'hf9b,
12'hfd5,
12'h013,
12'h009,
12'hf91,
12'hef1,
12'he8a,
12'he5a,
12'he5f,
12'heb8,
12'hf34,
12'hf8c,
12'hf81,
12'hf1f,
12'hed6,
12'hee1,
12'hf0e,
12'heff,
12'he95,
12'he1c,
12'hde3,
12'hde1,
12'he05,
12'he51,
12'heb5,
12'hef6,
12'hee5,
12'he9f,
12'he6d,
12'he85,
12'hecf,
12'hf11,
12'hf24,
12'hf1b,
12'hf03,
12'hedc,
12'hebb,
12'hec7,
12'hf09,
12'hf59,
12'hf7d,
12'hf6c,
12'hf55,
12'hf4c,
12'hf57,
12'hf66,
12'hf74,
12'hf90,
12'hf97,
12'hf78,
12'hf55,
12'hf6f,
12'hfd1,
12'h027,
12'h05e,
12'h08e,
12'h0c4,
12'h0eb,
12'h0da,
12'h0a6,
12'h0a5,
12'h101,
12'h167,
12'h192,
12'h17e,
12'h152,
12'h129,
12'h0fe,
12'h0e8,
12'h105,
12'h149,
12'h175,
12'h16d,
12'h128,
12'h0da,
12'h0ac,
12'h0aa,
12'h0d5,
12'h0fe,
12'h113,
12'h104,
12'h0e7,
12'h0c6,
12'h0af,
12'h0ac,
12'h0be,
12'h0c5,
12'h098,
12'h05a,
12'h023,
12'hffc,
12'hff2,
12'h012,
12'h049,
12'h058,
12'h00b,
12'hf9a,
12'hf54,
12'hf49,
12'hf4f,
12'hf40,
12'hf1d,
12'heef,
12'heaf,
12'he70,
12'he70,
12'hebb,
12'hf20,
12'hf49,
12'hf16,
12'hec4,
12'he79,
12'he42,
12'he37,
12'he49,
12'he73,
12'he93,
12'he83,
12'he74,
12'he84,
12'hed3,
12'hf4b,
12'hf99,
12'hf97,
12'hf50,
12'hee8,
12'he89,
12'he3e,
12'he10,
12'he1a,
12'he50,
12'he7d,
12'he7f,
12'he7e,
12'heb3,
12'hf14,
12'hf6a,
12'hfaa,
12'hfb6,
12'hf7a,
12'hf05,
12'he86,
12'he57,
12'he92,
12'hef9,
12'hf4e,
12'hf82,
12'hfaf,
12'hffb,
12'h067,
12'h0c1,
12'h0de,
12'h0bc,
12'h054,
12'hfc7,
12'hf61,
12'hf56,
12'hfa0,
12'hfff,
12'h05b,
12'h0b0,
12'h0fb,
12'h14c,
12'h1a9,
12'h200,
12'h224,
12'h208,
12'h1a9,
12'h11d,
12'h0c2,
12'h0f3,
12'h19a,
12'h24a,
12'h2b2,
12'h2ec,
12'h30f,
12'h311,
12'h308,
12'h2f6,
12'h2db,
12'h2a3,
12'h246,
12'h1ea,
12'h1a6,
12'h18f,
12'h1a6,
12'h1d5,
12'h1f4,
12'h1e4,
12'h1ac,
12'h170,
12'h15e,
12'h173,
12'h181,
12'h165,
12'h123,
12'h0c9,
12'h070,
12'h046,
12'h04d,
12'h072,
12'h095,
12'h099,
12'h081,
12'h053,
12'h023,
12'hfec,
12'hf9c,
12'hf36,
12'hed8,
12'heba,
12'hed8,
12'hf1b,
12'hf6b,
12'hfb0,
12'hfca,
12'hf96,
12'hf4b,
12'hf1e,
12'hf0c,
12'hefa,
12'heba,
12'he6c,
12'he49,
12'he48,
12'he68,
12'he9f,
12'hee1,
12'hf13,
12'hf02,
12'heb6,
12'he83,
12'hea4,
12'hefa,
12'hf4c,
12'hf72,
12'hf6e,
12'hf40,
12'hee1,
12'he8c,
12'hea5,
12'hf31,
12'hfc4,
12'h000,
12'hfe5,
12'hfa6,
12'hf74,
12'hf71,
12'hf8e,
12'hfae,
12'hfb4,
12'hf8b,
12'hf2c,
12'hed7,
12'hed2,
12'hf3b,
12'h004,
12'h0bf,
12'h102,
12'h0d1,
12'h066,
12'h00e,
12'h00e,
12'h06a,
12'h0f6,
12'h15b,
12'h157,
12'h103,
12'h0ae,
12'h091,
12'h0a5,
12'h0c9,
12'h0e6,
12'h0f7,
12'h0dc,
12'h090,
12'h04c,
12'h048,
12'h081,
12'h0ad,
12'h0a7,
12'h084,
12'h068,
12'h065,
12'h075,
12'h08a,
12'h098,
12'h091,
12'h07a,
12'h053,
12'h00b,
12'hfd3,
12'hfb8,
12'hfa5,
12'hf83,
12'hf67,
12'hf7e,
12'hfaf,
12'hfd1,
12'hfe0,
12'hfda,
12'hfb7,
12'hf66,
12'heee,
12'he99,
12'he84,
12'he89,
12'he8b,
12'he8a,
12'he9d,
12'hec0,
12'hee2,
12'heea,
12'hee4,
12'hed9,
12'hec1,
12'he8b,
12'he47,
12'he38,
12'he6e,
12'heb5,
12'hee7,
12'hefe,
12'hf12,
12'hf28,
12'hf2a,
12'hf37,
12'hf55,
12'hf7e,
12'hfa1,
12'hf8e,
12'hf32,
12'hed4,
12'heba,
12'hece,
12'heec,
12'hf17,
12'hf54,
12'hf75,
12'hf56,
12'hf16,
12'hf0f,
12'hf3b,
12'hf4f,
12'hf27,
12'hece,
12'he8e,
12'he92,
12'heef,
12'hf8b,
12'h047,
12'h0f3,
12'h14d,
12'h137,
12'h0c8,
12'h050,
12'hff9,
12'hfbb,
12'hf90,
12'hf70,
12'hf65,
12'hf7a,
12'hfbf,
12'h061,
12'h14d,
12'h229,
12'h29a,
12'h289,
12'h22e,
12'h1c8,
12'h172,
12'h128,
12'h0f8,
12'h103,
12'h152,
12'h1c0,
12'h224,
12'h283,
12'h2ef,
12'h34e,
12'h378,
12'h34f,
12'h2e8,
12'h28d,
12'h254,
12'h228,
12'h20b,
12'h1f5,
12'h1d0,
12'h1ab,
12'h197,
12'h192,
12'h19d,
12'h1c1,
12'h1eb,
12'h203,
12'h1ee,
12'h195,
12'h117,
12'h0a4,
12'h062,
12'h042,
12'h02b,
12'h020,
12'h018,
12'h010,
12'h016,
12'h026,
12'h045,
12'h04c,
12'h01f,
12'hfba,
12'hf2f,
12'hed4,
12'heb2,
12'hebd,
12'hefc,
12'hf59,
12'hf88,
12'hf46,
12'hede,
12'heaf,
12'hec3,
12'hedd,
12'heb6,
12'he7f,
12'he69,
12'he62,
12'he5a,
12'he5d,
12'he96,
12'heed,
12'hf23,
12'hf16,
12'hee4,
12'hecf,
12'hee9,
12'hf13,
12'hf32,
12'hf42,
12'hf2c,
12'hed7,
12'he6a,
12'he46,
12'he8c,
12'hf04,
12'hf6b,
12'hfab,
12'hfcb,
12'hfcc,
12'hfc8,
12'hfce,
12'hfd6,
12'hfd9,
12'hfbd,
12'hf71,
12'hf10,
12'hee4,
12'hf2c,
12'hfc6,
12'h053,
12'h0a8,
12'h0d8,
12'h0ec,
12'h0d6,
12'h0ab,
12'h0a1,
12'h0f1,
12'h167,
12'h195,
12'h167,
12'h126,
12'h10a,
12'h108,
12'h10b,
12'h125,
12'h15b,
12'h181,
12'h169,
12'h10d,
12'h0a8,
12'h07c,
12'h085,
12'h092,
12'h098,
12'h0a0,
12'h0a9,
12'h0c3,
12'h0dd,
12'h0ea,
12'h0f5,
12'h0f6,
12'h0e1,
12'h09e,
12'h044,
12'h002,
12'hfe1,
12'hfd9,
12'hfdb,
12'hfdc,
12'hfd3,
12'hfba,
12'hf96,
12'hf7d,
12'hf8a,
12'hf91,
12'hf6b,
12'hf24,
12'hed3,
12'he81,
12'he33,
12'he0c,
12'he24,
12'he7a,
12'hed7,
12'hefb,
12'hedd,
12'heb7,
12'heb1,
12'heb8,
12'heb4,
12'hea2,
12'heac,
12'hecf,
12'heea,
12'hee0,
12'hebb,
12'heb6,
12'hec8,
12'hed4,
12'hec7,
12'hea2,
12'he8c,
12'he7a,
12'he55,
12'he39,
12'he33,
12'he3e,
12'he59,
12'he7d,
12'heb8,
12'hf03,
12'hf51,
12'hf89,
12'hf98,
12'hf94,
12'hf7c,
12'hf43,
12'hee9,
12'hea2,
12'he8d,
12'hea6,
12'heee,
12'hf50,
12'hfd5,
12'h060,
12'h0b6,
12'h0bf,
12'h084,
12'h032,
12'hfdc,
12'hf94,
12'hf69,
12'hf62,
12'hf82,
12'hfb0,
12'hfdb,
12'h02b,
12'h0cc,
12'h179,
12'h1eb,
12'h21d,
12'h23b,
12'h25b,
12'h249,
12'h209,
12'h1e3,
12'h1fd,
12'h236,
12'h24c,
12'h25e,
12'h2a7,
12'h306,
12'h33b,
12'h322,
12'h2dd,
12'h29f,
12'h270,
12'h24f,
12'h24d,
12'h24c,
12'h236,
12'h206,
12'h1ce,
12'h1ac,
12'h18f,
12'h181,
12'h18d,
12'h1a9,
12'h1b6,
12'h196,
12'h163,
12'h12f,
12'h0fe,
12'h0d2,
12'h0ad,
12'h094,
12'h077,
12'h04d,
12'h02b,
12'h011,
12'h000,
12'hfe2,
12'hf8f,
12'hf22,
12'hed7,
12'heda,
12'hf09,
12'hf26,
12'hf4a,
12'hf85,
12'hfc1,
12'hfba,
12'hf65,
12'hf1a,
12'hefd,
12'heeb,
12'heb0,
12'he5f,
12'he3a,
12'he51,
12'he7f,
12'he9e,
12'head,
12'hebc,
12'heb6,
12'he96,
12'he81,
12'he9d,
12'heee,
12'hf3c,
12'hf68,
12'hf80,
12'hf76,
12'hf43,
12'hf01,
12'heec,
12'hf16,
12'hf49,
12'hf4e,
12'hf31,
12'hf24,
12'hf43,
12'hf85,
12'hfc9,
12'hffc,
12'h01e,
12'h020,
12'hfe9,
12'hf93,
12'hf64,
12'hf91,
12'h005,
12'h062,
12'h085,
12'h08c,
12'h098,
12'h09e,
12'h095,
12'h0b2,
12'h0fd,
12'h143,
12'h155,
12'h13f,
12'h126,
12'h10e,
12'h0f3,
12'h0df,
12'h0ef,
12'h117,
12'h122,
12'h100,
12'h0c4,
12'h096,
12'h093,
12'h0aa,
12'h0c5,
12'h0cb,
12'h0b9,
12'h0a1,
12'h086,
12'h068,
12'h056,
12'h060,
12'h069,
12'h059,
12'h03a,
12'h00a,
12'hfdd,
12'hfc6,
12'hfbb,
12'hfaf,
12'hf9f,
12'hf88,
12'hf67,
12'hf3e,
12'hf22,
12'hf22,
12'hf24,
12'hf06,
12'hecc,
12'hea5,
12'he92,
12'he73,
12'he49,
12'he3d,
12'he6f,
12'hea6,
12'head,
12'he92,
12'he81,
12'he81,
12'he80,
12'he76,
12'he5c,
12'he5b,
12'he86,
12'hecc,
12'hf06,
12'hf2a,
12'hf56,
12'hf79,
12'hf8c,
12'hf9a,
12'hf9e,
12'hf7b,
12'hf1b,
12'hea5,
12'he62,
12'he71,
12'hec1,
12'hf21,
12'hf5e,
12'hf60,
12'hf34,
12'hf04,
12'hef9,
12'hf1b,
12'hf46,
12'hf4a,
12'hf0f,
12'hebb,
12'hea3,
12'hef7,
12'hf84,
12'h002,
12'h06d,
12'h0d2,
12'h105,
12'h0de,
12'h090,
12'h058,
12'h044,
12'h028,
12'hfe8,
12'hfaf,
12'hfab,
12'hfe6,
12'h044,
12'h0c3,
12'h150,
12'h1b8,
12'h1d6,
12'h1b6,
12'h18a,
12'h17b,
12'h18d,
12'h19a,
12'h192,
12'h190,
12'h1c9,
12'h23e,
12'h2bf,
12'h33f,
12'h3a0,
12'h3c3,
12'h39c,
12'h330,
12'h2ad,
12'h233,
12'h1d5,
12'h1a5,
12'h19d,
12'h19a,
12'h196,
12'h1ae,
12'h1dd,
12'h20c,
12'h221,
12'h212,
12'h1e8,
12'h196,
12'h11c,
12'h099,
12'h03d,
12'h019,
12'h021,
12'h042,
12'h06f,
12'h080,
12'h07b,
12'h077,
12'h06f,
12'h061,
12'h030,
12'hfda,
12'hf5b,
12'hecf,
12'he69,
12'he30,
12'he32,
12'he65,
12'hebb,
12'hf0f,
12'hf2e,
12'hf12,
12'hee5,
12'heee,
12'hf14,
12'hf1f,
12'heea,
12'he7e,
12'he2d,
12'he06,
12'hdff,
12'he24,
12'he73,
12'hec6,
12'heeb,
12'hedc,
12'hed4,
12'hef2,
12'hf20,
12'hf49,
12'hf56,
12'hf45,
12'hf0e,
12'heae,
12'he5a,
12'he56,
12'hebb,
12'hf48,
12'hfac,
12'hfd4,
12'hfd4,
12'hfbe,
12'hfa3,
12'hfa2,
12'hfaf,
12'hfc0,
12'hfc1,
12'hf90,
12'hf4f,
12'hf44,
12'hf98,
12'h01d,
12'h099,
12'h0f1,
12'h116,
12'h10f,
12'h0d4,
12'h091,
12'h08f,
12'h0dc,
12'h13b,
12'h166,
12'h154,
12'h12b,
12'h111,
12'h10a,
12'h11e,
12'h155,
12'h192,
12'h1b1,
12'h18a,
12'h122,
12'h0b8,
12'h090,
12'h0a3,
12'h0bc,
12'h0c5,
12'h0c5,
12'h0c9,
12'h0c9,
12'h0ca,
12'h0db,
12'h0ff,
12'h114,
12'h0f7,
12'h0ae,
12'h055,
12'h019,
12'h000,
12'hff5,
12'hffc,
12'h010,
12'h016,
12'hffa,
12'hfca,
12'hfa7,
12'hf9c,
12'hf88,
12'hf3c,
12'hec9,
12'he68,
12'he2a,
12'he00,
12'hdf0,
12'he22,
12'he85,
12'hed4,
12'hee4,
12'hec4,
12'heba,
12'hecd,
12'hecb,
12'hea1,
12'he70,
12'he68,
12'he77,
12'he6e,
12'he54,
12'he63,
12'heaf,
12'hf03,
12'hf20,
12'hf20,
12'hf27,
12'hf25,
12'hf05,
12'heab,
12'he4f,
12'he24,
12'he33,
12'he6f,
12'hebc,
12'hf07,
12'hf3f,
12'hf74,
12'hfa3,
12'hfd4,
12'h000,
12'hff1,
12'hf85,
12'hedc,
12'he6a,
12'he67,
12'heb2,
12'hf1d,
12'hf7b,
12'hfd6,
12'h026,
12'h068,
12'h0a6,
12'h0e2,
12'h0fb,
12'h0c9,
12'h050,
12'hfc0,
12'hf6d,
12'hf78,
12'hfc0,
12'h029,
12'h0a5,
12'h12c,
12'h193,
12'h1bf,
12'h1c7,
12'h1e2,
12'h232,
12'h254,
12'h21b,
12'h1cf,
12'h1c2,
12'h200,
12'h245,
12'h27e,
12'h2c0,
12'h2f6,
12'h2e9,
12'h2a6,
12'h275,
12'h26f,
12'h27e,
12'h28b,
12'h276,
12'h22a,
12'h1ca,
12'h18c,
12'h17b,
12'h17a,
12'h165,
12'h145,
12'h132,
12'h12c,
12'h125,
12'h11a,
12'h112,
12'h0ff,
12'h0da,
12'h0a6,
12'h071,
12'h042,
12'h017,
12'hff3,
12'hfdb,
12'hfc5,
12'hf99,
12'hf52,
12'hf01,
12'hec5,
12'heb4,
12'hecf,
12'hefe,
12'hf28,
12'hf56,
12'hf7b,
12'hf76,
12'hf32,
12'heda,
12'heaa,
12'he9c,
12'he90,
12'he63,
12'he2c,
12'he2a,
12'he54,
12'he7b,
12'he94,
12'hebf,
12'hef8,
12'hf0c,
12'hed0,
12'he75,
12'he66,
12'heab,
12'hf0e,
12'hf4c,
12'hf5c,
12'hf46,
12'hf08,
12'hebc,
12'he95,
12'hed1,
12'hf3c,
12'hf8d,
12'hfa6,
12'hf97,
12'hf8d,
12'hf95,
12'hfbd,
12'hffa,
12'h033,
12'h047,
12'h006,
12'hf98,
12'hf61,
12'hf9a,
12'h017,
12'h083,
12'h0bb,
12'h0cc,
12'h0b9,
12'h07f,
12'h052,
12'h081,
12'h11e,
12'h1c2,
12'h1e8,
12'h18c,
12'h117,
12'h0d9,
12'h0de,
12'h104,
12'h135,
12'h166,
12'h176,
12'h148,
12'h0f0,
12'h0b6,
12'h0d1,
12'h11e,
12'h146,
12'h11c,
12'h0c4,
12'h07b,
12'h05f,
12'h072,
12'h094,
12'h0ae,
12'h0bf,
12'h0b8,
12'h088,
12'h03c,
12'h00b,
12'h00a,
12'h01c,
12'h024,
12'h005,
12'hfd1,
12'hf98,
12'hf62,
12'hf4b,
12'hf51,
12'hf52,
12'hf28,
12'hed4,
12'he8d,
12'he72,
12'he64,
12'he6d,
12'hea6,
12'hef0,
12'hf04,
12'hec7,
12'he78,
12'he56,
12'he6b,
12'he7e,
12'he67,
12'he4e,
12'he64,
12'he99,
12'heb5,
12'heb5,
12'hec0,
12'hed9,
12'hed5,
12'he98,
12'he4d,
12'he25,
12'he27,
12'he41,
12'he53,
12'he63,
12'he92,
12'hee5,
12'hf32,
12'hf6a,
12'hfab,
12'hff9,
12'h036,
12'h027,
12'hfc4,
12'hf47,
12'hed9,
12'he7e,
12'he38,
12'he20,
12'he49,
12'he97,
12'hee8,
12'hf39,
12'hfb7,
12'h06a,
12'h115,
12'h168,
12'h149,
12'h0c6,
12'h010,
12'hf6e,
12'hf14,
12'hf1e,
12'hf6c,
12'hfcc,
12'h02d,
12'h0aa,
12'h156,
12'h211,
12'h29e,
12'h2db,
12'h2c9,
12'h263,
12'h1c0,
12'h11b,
12'h0c0,
12'h0f2,
12'h185,
12'h1fa,
12'h232,
12'h25d,
12'h29d,
12'h2e3,
12'h310,
12'h321,
12'h30c,
12'h2c2,
12'h258,
12'h1fb,
12'h1c3,
12'h1a9,
12'h1ad,
12'h1bb,
12'h1b7,
12'h196,
12'h16b,
12'h164,
12'h196,
12'h1db,
12'h1ea,
12'h1a0,
12'h11c,
12'h08d,
12'h023,
12'hff6,
12'hfee,
12'hff2,
12'hfef,
12'hfd8,
12'hfbd,
12'hfb1,
12'hfb8,
12'hfc5,
12'hfb1,
12'hf66,
12'hf0c,
12'hec8,
12'hebc,
12'hef3,
12'hf53,
12'hfa2,
12'hf9a,
12'hf49,
12'hef3,
12'hecf,
12'hed5,
12'hec8,
12'he9c,
12'he71,
12'he5e,
12'he50,
12'he42,
12'he50,
12'he90,
12'hedc,
12'hef2,
12'hed6,
12'hec8,
12'hefd,
12'hf5b,
12'hfa2,
12'hfbb,
12'hfab,
12'hf7e,
12'hf25,
12'hec5,
12'heb3,
12'hef8,
12'hf5c,
12'hfa5,
12'hfc2,
12'hfc4,
12'hfc3,
12'hfd6,
12'h001,
12'h035,
12'h04b,
12'h019,
12'hfb0,
12'hf5d,
12'hf6d,
12'hfdb,
12'h05e,
12'h0b3,
12'h0cb,
12'h0c1,
12'h0ae,
12'h0a3,
12'h0bd,
12'h10d,
12'h166,
12'h185,
12'h14e,
12'h0f9,
12'h0d1,
12'h0e8,
12'h114,
12'h130,
12'h149,
12'h163,
12'h170,
12'h160,
12'h13d,
12'h121,
12'h107,
12'h0db,
12'h09a,
12'h05f,
12'h040,
12'h053,
12'h07c,
12'h090,
12'h096,
12'h0a2,
12'h0be,
12'h0d1,
12'h0bf,
12'h08f,
12'h04b,
12'hff3,
12'hf96,
12'hf5e,
12'hf66,
12'hf84,
12'hf6e,
12'hf35,
12'hf1a,
12'hf2a,
12'hf3d,
12'hf30,
12'hf18,
12'hf0c,
12'heed,
12'hea1,
12'he4f,
12'he31,
12'he4b,
12'he67,
12'he55,
12'he31,
12'he21,
12'he29,
12'he33,
12'he34,
12'he5d,
12'heb6,
12'hf00,
12'hf15,
12'hef5,
12'hecb,
12'heaf,
12'he96,
12'he8e,
12'he98,
12'hea7,
12'heb0,
12'heab,
12'heab,
12'hec4,
12'hee4,
12'hee9,
12'hecd,
12'hecc,
12'hef8,
12'hf33,
12'hf50,
12'hf3e,
12'hf1e,
12'heff,
12'hee8,
12'hedf,
12'hef4,
12'hf20,
12'hf47,
12'hf69,
12'hf87,
12'hfc7,
12'h039,
12'h09c,
12'h0c0,
12'h0a0,
12'h059,
12'h00e,
12'hfdf,
12'hfe3,
12'h01e,
12'h075,
12'h0a9,
12'h09d,
12'h0a3,
12'h0fe,
12'h183,
12'h1e7,
12'h203,
12'h1ee,
12'h1d7,
12'h1b6,
12'h190,
12'h198,
12'h1f2,
12'h289,
12'h301,
12'h31c,
12'h314,
12'h31b,
12'h32d,
12'h321,
12'h2d6,
12'h280,
12'h23c,
12'h201,
12'h1ec,
12'h204,
12'h239,
12'h264,
12'h268,
12'h25d,
12'h245,
12'h208,
12'h1b3,
12'h16f,
12'h151,
12'h139,
12'h0fe,
12'h0ae,
12'h073,
12'h070,
12'h090,
12'h0a4,
12'h0a0,
12'h09c,
12'h093,
12'h077,
12'h04f,
12'h01a,
12'hfcd,
12'hf4b,
12'heb1,
12'he5e,
12'he69,
12'he99,
12'hec4,
12'hefc,
12'hf46,
12'hf6b,
12'hf56,
12'hf45,
12'hf4d,
12'hf49,
12'hefd,
12'he68,
12'hdf8,
12'hde8,
12'he1a,
12'he5e,
12'he8d,
12'heb5,
12'heeb,
12'hefe,
12'hed9,
12'hec3,
12'hedb,
12'heff,
12'hf0f,
12'hf08,
12'hf01,
12'heef,
12'heca,
12'heb0,
12'hedf,
12'hf3b,
12'hf6c,
12'hf6c,
12'hf52,
12'hf4c,
12'hf75,
12'hfac,
12'hfd4,
12'hfea,
12'hfed,
12'hfca,
12'hf75,
12'hf32,
12'hf4f,
12'hfc4,
12'h03a,
12'h068,
12'h052,
12'h039,
12'h036,
12'h04b,
12'h081,
12'h0d4,
12'h12c,
12'h153,
12'h132,
12'h0f2,
12'h0ce,
12'h0dc,
12'h0f2,
12'h0f9,
12'h0f8,
12'h0fc,
12'h103,
12'h0ef,
12'h0c8,
12'h0b7,
12'h0b8,
12'h0ad,
12'h094,
12'h085,
12'h08f,
12'h0aa,
12'h0be,
12'h0c1,
12'h0cd,
12'h0d4,
12'h0ba,
12'h07b,
12'h021,
12'hfe3,
12'hfcd,
12'hfc5,
12'hfc1,
12'hfbc,
12'hfc8,
12'hfd5,
12'hfb6,
12'hf80,
12'hf53,
12'hf28,
12'hee8,
12'heaa,
12'he98,
12'hea3,
12'hea3,
12'he8c,
12'he71,
12'he72,
12'he95,
12'hea8,
12'he90,
12'he74,
12'he77,
12'he8c,
12'he85,
12'he61,
12'he53,
12'he76,
12'hea0,
12'hea6,
12'he9c,
12'heb2,
12'heef,
12'hf37,
12'hf71,
12'hf77,
12'hf4d,
12'hf0e,
12'hec8,
12'he8c,
12'he5a,
12'he43,
12'he43,
12'he65,
12'hebc,
12'hf3d,
12'hfc4,
12'h018,
12'h01e,
12'hff8,
12'hfbd,
12'hf6d,
12'hf26,
12'heef,
12'hed2,
12'hedc,
12'hf05,
12'hf4b,
12'hfbc,
12'h04c,
12'h0c6,
12'h0f5,
12'h0cf,
12'h08a,
12'h04c,
12'h01b,
12'hffd,
12'hff4,
12'h016,
12'h039,
12'h03c,
12'h062,
12'h0d9,
12'h184,
12'h212,
12'h24f,
12'h24d,
12'h232,
12'h217,
12'h1ee,
12'h1d8,
12'h204,
12'h258,
12'h295,
12'h292,
12'h28a,
12'h2b9,
12'h308,
12'h33a,
12'h32b,
12'h2f4,
12'h290,
12'h200,
12'h19c,
12'h19f,
12'h1ee,
12'h22b,
12'h221,
12'h203,
12'h1ec,
12'h1cc,
12'h1af,
12'h1a9,
12'h1b1,
12'h19e,
12'h147,
12'h0c9,
12'h064,
12'h03d,
12'h04d,
12'h067,
12'h070,
12'h05e,
12'h036,
12'h007,
12'hfff,
12'h018,
12'h00d,
12'hfb9,
12'hf1b,
12'he85,
12'he42,
12'he44,
12'he76,
12'hedf,
12'hf64,
12'hf9e,
12'hf69,
12'hf02,
12'hebc,
12'hec0,
12'hecf,
12'hea8,
12'he62,
12'he47,
12'he57,
12'he6f,
12'he8c,
12'heac,
12'hed1,
12'hed7,
12'hea8,
12'he70,
12'he62,
12'he8d,
12'hed9,
12'hf30,
12'hf62,
12'hf4f,
12'hef5,
12'he96,
12'he85,
12'hec1,
12'hf1e,
12'hf65,
12'hf86,
12'hf9c,
12'hfb1,
12'hfd6,
12'hff2,
12'hff5,
12'hfeb,
12'hfcc,
12'hf8f,
12'hf48,
12'hf43,
12'hf9e,
12'h01f,
12'h081,
12'h0ad,
12'h0c8,
12'h0dc,
12'h0cc,
12'h09b,
12'h086,
12'h0c9,
12'h136,
12'h17b,
12'h176,
12'h143,
12'h10b,
12'h0d7,
12'h0b5,
12'h0c6,
12'h10b,
12'h14e,
12'h156,
12'h11d,
12'h0d4,
12'h0a7,
12'h099,
12'h0ac,
12'h0cf,
12'h0e7,
12'h0e5,
12'h0c8,
12'h0ab,
12'h0ab,
12'h0bf,
12'h0cd,
12'h0bc,
12'h07e,
12'h02e,
12'hff3,
12'hfd0,
12'hfc6,
12'hfc7,
12'hfdf,
12'h008,
12'h014,
12'hfe2,
12'hf82,
12'hf35,
12'hf0d,
12'hef6,
12'hee9,
12'hee0,
12'hec8,
12'he97,
12'he67,
12'he63,
12'he9b,
12'heec,
12'hf0a,
12'heeb,
12'heb7,
12'he89,
12'he74,
12'he5f,
12'he51,
12'he68,
12'he8b,
12'he91,
12'he7e,
12'he8a,
12'hed2,
12'hf36,
12'hf85,
12'hfa2,
12'hf87,
12'hf3b,
12'hed7,
12'he6b,
12'he2b,
12'he4b,
12'hea3,
12'hee1,
12'hee5,
12'hedc,
12'hf0b,
12'hf62,
12'hfa3,
12'hfb3,
12'hfa0,
12'hf5f,
12'hef0,
12'he8c,
12'he78,
12'hec8,
12'hf46,
12'hfa9,
12'hfe5,
12'h01f,
12'h061,
12'h08e,
12'h099,
12'h094,
12'h076,
12'h025,
12'hfc8,
12'hfa1,
12'hfca,
12'h010,
12'h046,
12'h08a,
12'h0f9,
12'h171,
12'h1c3,
12'h1da,
12'h1ce,
12'h1c0,
12'h191,
12'h14f,
12'h12c,
12'h149,
12'h1b6,
12'h23e,
12'h2a1,
12'h2d6,
12'h303,
12'h333,
12'h34f,
12'h345,
12'h30a,
12'h29b,
12'h20b,
12'h195,
12'h155,
12'h144,
12'h166,
12'h1a1,
12'h1de,
12'h1f8,
12'h1d1,
12'h1aa,
12'h1ab,
12'h1b8,
12'h19c,
12'h143,
12'h0d4,
12'h06b,
12'h01e,
12'hff5,
12'hfff,
12'h021,
12'h02d,
12'h02c,
12'h02d,
12'h03c,
12'h047,
12'h037,
12'h001,
12'hf8e,
12'hefd,
12'he91,
12'he68,
12'he88,
12'hed3,
12'hf20,
12'hf3e,
12'hf17,
12'hee7,
12'heed,
12'hf12,
12'hf2a,
12'hf1c,
12'hee9,
12'heab,
12'he7d,
12'he69,
12'he77,
12'heaa,
12'hee3,
12'hef5,
12'hed5,
12'hea4,
12'he9d,
12'hee8,
12'hf57,
12'hf9f,
12'hfad,
12'hf86,
12'hf26,
12'hebc,
12'he95,
12'hed8,
12'hf5c,
12'hfc7,
12'hfe0,
12'hfb7,
12'hf96,
12'hfab,
12'hfd7,
12'hfeb,
12'hfe2,
12'hfc9,
12'hfa1,
12'hf6c,
12'hf57,
12'hf98,
12'h018,
12'h09f,
12'h0eb,
12'h0f7,
12'h0d2,
12'h08d,
12'h04d,
12'h049,
12'h0a7,
12'h121,
12'h168,
12'h15d,
12'h11e,
12'h0f5,
12'h0f2,
12'h0ff,
12'h118,
12'h136,
12'h14e,
12'h13a,
12'h0ec,
12'h0a4,
12'h089,
12'h098,
12'h0ad,
12'h0ad,
12'h0a0,
12'h09c,
12'h0ae,
12'h0bf,
12'h0be,
12'h0b5,
12'h0be,
12'h0c7,
12'h097,
12'h02f,
12'hfcc,
12'hf8f,
12'hf86,
12'hf98,
12'hfbd,
12'hff0,
12'hffe,
12'hfd6,
12'hfa2,
12'hf7e,
12'hf57,
12'hf11,
12'hec1,
12'he92,
12'he73,
12'he4d,
12'he20,
12'he0e,
12'he40,
12'he88,
12'hea7,
12'he92,
12'he7a,
12'he90,
12'heb1,
12'heab,
12'he8e,
12'he88,
12'he9d,
12'heab,
12'hea4,
12'he93,
12'he93,
12'hec2,
12'hefe,
12'hf30,
12'hf41,
12'hf2f,
12'hf15,
12'hee7,
12'heac,
12'he74,
12'he5e,
12'he62,
12'he78,
12'heb6,
12'hf17,
12'hf82,
12'hfc6,
12'hfdb,
12'hfd1,
12'hfb7,
12'hf94,
12'hf61,
12'hf1d,
12'hee0,
12'hece,
12'hef0,
12'hf41,
12'hfae,
12'h028,
12'h096,
12'h0c7,
12'h0be,
12'h0ac,
12'h09c,
12'h07c,
12'h046,
12'h00c,
12'hff7,
12'h00d,
12'h03a,
12'h089,
12'h109,
12'h194,
12'h1e5,
12'h1d8,
12'h1ae,
12'h1be,
12'h1ff,
12'h221,
12'h209,
12'h201,
12'h234,
12'h276,
12'h2a8,
12'h2e3,
12'h32b,
12'h349,
12'h310,
12'h291,
12'h222,
12'h1ec,
12'h1e2,
12'h200,
12'h224,
12'h229,
12'h1f8,
12'h1ba,
12'h1a8,
12'h1b4,
12'h1b8,
12'h19f,
12'h170,
12'h134,
12'h0f0,
12'h0b4,
12'h094,
12'h092,
12'h095,
12'h080,
12'h04d,
12'h018,
12'hffc,
12'hffc,
12'h003,
12'h004,
12'hfe4,
12'hf84,
12'heed,
12'he59,
12'he31,
12'he77,
12'hec7,
12'hefb,
12'hf24,
12'hf53,
12'hf62,
12'hf3c,
12'hf11,
12'hf05,
12'hf06,
12'hecd,
12'he4f,
12'hdea,
12'hde7,
12'he28,
12'he64,
12'he8b,
12'heb3,
12'hedf,
12'hee2,
12'hebb,
12'hea5,
12'hecc,
12'hf09,
12'hf25,
12'hf2e,
12'hf36,
12'hf39,
12'hf0b,
12'hec4,
12'hec1,
12'hf05,
12'hf4b,
12'hf73,
12'hf90,
12'hfad,
12'hfba,
12'hfbe,
12'hfc2,
12'hfd1,
12'hff2,
12'hffe,
12'hfd7,
12'hf8f,
12'hf70,
12'hfab,
12'h01c,
12'h07a,
12'h0a7,
12'h0c1,
12'h0c0,
12'h096,
12'h062,
12'h075,
12'h0fa,
12'h190,
12'h1d1,
12'h19f,
12'h13b,
12'h0f3,
12'h0db,
12'h0f2,
12'h12a,
12'h173,
12'h18f,
12'h155,
12'h0e5,
12'h091,
12'h08d,
12'h0c1,
12'h0ef,
12'h0fc,
12'h0e7,
12'h0bb,
12'h09f,
12'h0a5,
12'h0c9,
12'h0ed,
12'h0f0,
12'h0bb,
12'h04f,
12'hfe5,
12'hfb7,
12'hfd2,
12'h007,
12'h031,
12'h039,
12'h019,
12'hfd6,
12'hf74,
12'hf38,
12'hf3a,
12'hf46,
12'hf1e,
12'hebf,
12'he70,
12'he4c,
12'he4c,
12'he54,
12'he6b,
12'hea2,
12'hed3,
12'hed0,
12'hea7,
12'he96,
12'heae,
12'hebe,
12'he93,
12'he45,
12'he18,
12'he2d,
12'he52,
12'he78,
12'heb4,
12'hf09,
12'hf58,
12'hf8a,
12'hf88,
12'hf5b,
12'hf26,
12'hee3,
12'he8d,
12'he3c,
12'he28,
12'he45,
12'he67,
12'he97,
12'hefe,
12'hf98,
12'h00a,
12'h011,
12'hfdc,
12'hf99,
12'hf42,
12'hee7,
12'heb0,
12'heb4,
12'hed6,
12'hefa,
12'hf1d,
12'hf61,
12'hfd8,
12'h060,
12'h0cc,
12'h0f2,
12'h0cc,
12'h071,
12'h012,
12'hfe6,
12'hfe7,
12'hff6,
12'hffd,
12'h003,
12'h034,
12'h097,
12'h123,
12'h1b7,
12'h218,
12'h229,
12'h1fa,
12'h1c5,
12'h1b9,
12'h1ce,
12'h1f0,
12'h22a,
12'h268,
12'h279,
12'h267,
12'h27a,
12'h2da,
12'h340,
12'h359,
12'h318,
12'h2ab,
12'h249,
12'h20d,
12'h201,
12'h214,
12'h21e,
12'h200,
12'h1c7,
12'h188,
12'h15e,
12'h170,
12'h1b1,
12'h1de,
12'h1c8,
12'h176,
12'h110,
12'h0ba,
12'h083,
12'h073,
12'h075,
12'h066,
12'h02e,
12'hfea,
12'hfcf,
12'hfde,
12'hffd,
12'h002,
12'hfc5,
12'hf37,
12'he96,
12'he4f,
12'he7e,
12'hedb,
12'hf2f,
12'hf64,
12'hf69,
12'hf35,
12'hee0,
12'heb3,
12'hec8,
12'hef6,
12'hee6,
12'he82,
12'he1d,
12'hdfc,
12'he1d,
12'he5d,
12'hea2,
12'hed9,
12'hee4,
12'heaa,
12'he58,
12'he4c,
12'head,
12'hf2d,
12'hf6d,
12'hf78,
12'hf5e,
12'hf07,
12'he8f,
12'he53,
12'he92,
12'hf17,
12'hf7a,
12'hf92,
12'hf84,
12'hf83,
12'hf9b,
12'hfb5,
12'hfc3,
12'hfc0,
12'hfb1,
12'hf95,
12'hf65,
12'hf4b,
12'hf77,
12'hff4,
12'h076,
12'h0c0,
12'h0ca,
12'h0b6,
12'h09f,
12'h07c,
12'h071,
12'h0a3,
12'h0f0,
12'h13c,
12'h160,
12'h14d,
12'h12d,
12'h114,
12'h104,
12'h0fc,
12'h115,
12'h15d,
12'h196,
12'h17c,
12'h120,
12'h0cc,
12'h0a7,
12'h0a3,
12'h0a9,
12'h0c1,
12'h0db,
12'h0d2,
12'h0ad,
12'h08b,
12'h09a,
12'h0d8,
12'h0ff,
12'h0d8,
12'h072,
12'h005,
12'hfba,
12'hfa5,
12'hfb8,
12'hfe0,
12'h004,
12'hff5,
12'hfaf,
12'hf5b,
12'hf33,
12'hf34,
12'hf29,
12'hf0c,
12'hedf,
12'heac,
12'he69,
12'he2a,
12'he10,
12'he35,
12'he89,
12'hec5,
12'hec9,
12'hea0,
12'he8f,
12'he98,
12'he88,
12'he6a,
12'he59,
12'he67,
12'he7e,
12'he7e,
12'he80,
12'heb0,
12'hf0f,
12'hf65,
12'hf78,
12'hf4f,
12'hf0d,
12'hed5,
12'hea3,
12'he5c,
12'he1f,
12'he13,
12'he30,
12'he72,
12'hee0,
12'hf6c,
12'hfe3,
12'h00c,
12'hfee,
12'hfb4,
12'hf88,
12'hf60,
12'hf1b,
12'hed5,
12'heb9,
12'hede,
12'hf1e,
12'hf5c,
12'hfb9,
12'h043,
12'h0b9,
12'h0dd,
12'h0c8,
12'h0a2,
12'h072,
12'h02e,
12'hfe3,
12'hfbb,
12'hfd5,
12'h00b,
12'h047,
12'h0a3,
12'h132,
12'h1c8,
12'h233,
12'h25d,
12'h261,
12'h26b,
12'h24d,
12'h1eb,
12'h18c,
12'h186,
12'h1e3,
12'h259,
12'h2a5,
12'h2e4,
12'h328,
12'h349,
12'h32f,
12'h2ee,
12'h2b2,
12'h27b,
12'h244,
12'h220,
12'h209,
12'h1f6,
12'h1de,
12'h1c1,
12'h1bc,
12'h1af,
12'h17e,
12'h144,
12'h133,
12'h150,
12'h167,
12'h15a,
12'h11c,
12'h0cd,
12'h085,
12'h048,
12'h023,
12'h013,
12'h011,
12'h000,
12'hfdc,
12'hfbd,
12'hf93,
12'hf49,
12'hee7,
12'hea4,
12'hea3,
12'heae,
12'heac,
12'hec2,
12'hefa,
12'hf3a,
12'hf45,
12'hf14,
12'hee3,
12'hec9,
12'heb1,
12'he7c,
12'he3d,
12'he30,
12'he54,
12'he85,
12'heab,
12'heb9,
12'hec5,
12'hece,
12'heb5,
12'he7e,
12'he53,
12'he64,
12'hea3,
12'heea,
12'hf23,
12'hf44,
12'hf3a,
12'hf05,
12'hed6,
12'heda,
12'hf14,
12'hf54,
12'hf6d,
12'hf63,
12'hf58,
12'hf6d,
12'hf9c,
12'hfc9,
12'hfdd,
12'hfd4,
12'hfb2,
12'hf73,
12'hf47,
12'hf74,
12'hff4,
12'h07c,
12'h0af,
12'h09b,
12'h07f,
12'h075,
12'h066,
12'h060,
12'h0a4,
12'h12b,
12'h19d,
12'h1af,
12'h179,
12'h13e,
12'h11e,
12'h117,
12'h11d,
12'h138,
12'h15c,
12'h156,
12'h11a,
12'h0e5,
12'h0e8,
12'h10b,
12'h123,
12'h126,
12'h112,
12'h0e1,
12'h0b1,
12'h0b5,
12'h0e6,
12'h10d,
12'h10d,
12'h0ea,
12'h0a6,
12'h057,
12'h025,
12'h024,
12'h03c,
12'h03b,
12'h01e,
12'h009,
12'hffe,
12'hfdc,
12'hfa2,
12'hf6e,
12'hf4c,
12'hf2a,
12'hef5,
12'hec5,
12'heb2,
12'hea9,
12'he8e,
12'he70,
12'he7a,
12'heaa,
12'hed0,
12'hec6,
12'hea2,
12'he81,
12'he65,
12'he38,
12'hdff,
12'hdf3,
12'he2e,
12'he7d,
12'heac,
12'hebe,
12'hed9,
12'hf15,
12'hf51,
12'hf6c,
12'hf59,
12'hf24,
12'hed6,
12'he6b,
12'he0d,
12'hdfa,
12'he45,
12'hea6,
12'hecf,
12'hece,
12'hedf,
12'hf11,
12'hf53,
12'hf80,
12'hf77,
12'hf3a,
12'hee5,
12'he94,
12'he74,
12'head,
12'hf1c,
12'hf8a,
12'hfd4,
12'h00e,
12'h059,
12'h09a,
12'h0b2,
12'h09b,
12'h06b,
12'h01a,
12'hfa9,
12'hf54,
12'hf4f,
12'hf8b,
12'hfe5,
12'h04d,
12'h0d2,
12'h172,
12'h1fc,
12'h23d,
12'h23d,
12'h220,
12'h203,
12'h1d2,
12'h17e,
12'h130,
12'h12c,
12'h198,
12'h234,
12'h2b1,
12'h30b,
12'h34f,
12'h379,
12'h37a,
12'h344,
12'h2e4,
12'h279,
12'h21f,
12'h1dd,
12'h1a8,
12'h18c,
12'h1a1,
12'h1d8,
12'h20a,
12'h21a,
12'h202,
12'h1d9,
12'h1b9,
12'h1a4,
12'h181,
12'h14b,
12'h10c,
12'h0bb,
12'h072,
12'h04c,
12'h03c,
12'h034,
12'h03a,
12'h04c,
12'h054,
12'h04c,
12'h02f,
12'h001,
12'hfc4,
12'hf63,
12'hef3,
12'head,
12'hea6,
12'hec0,
12'hef3,
12'hf2b,
12'hf43,
12'hf35,
12'hf14,
12'hf10,
12'hf24,
12'hf0f,
12'hebb,
12'he62,
12'he2d,
12'he1c,
12'he36,
12'he81,
12'hede,
12'hf11,
12'hf05,
12'hecb,
12'he99,
12'hea0,
12'hed6,
12'hf0a,
12'hf19,
12'hf07,
12'hed8,
12'he90,
12'he56,
12'he68,
12'hed9,
12'hf6d,
12'hfce,
12'hfdf,
12'hfbe,
12'hf91,
12'hf7c,
12'hf8d,
12'hfbf,
12'hfe5,
12'hfdb,
12'hf99,
12'hf3c,
12'hf1b,
12'hf5e,
12'hfed,
12'h07a,
12'h0d2,
12'h0e4,
12'h0bc,
12'h07e,
12'h05d,
12'h087,
12'h0f8,
12'h165,
12'h183,
12'h153,
12'h107,
12'h0e5,
12'h102,
12'h13b,
12'h164,
12'h17e,
12'h175,
12'h135,
12'h0d4,
12'h08f,
12'h08c,
12'h0ac,
12'h0d4,
12'h0e3,
12'h0e0,
12'h0e3,
12'h0e8,
12'h0e9,
12'h0e2,
12'h0df,
12'h0d8,
12'h0b3,
12'h05e,
12'h003,
12'hfdc,
12'hfe7,
12'hff4,
12'hff1,
12'hfef,
12'hfe7,
12'hfc0,
12'hf8e,
12'hf73,
12'hf61,
12'hf35,
12'heed,
12'he9f,
12'he67,
12'he4a,
12'he2d,
12'he14,
12'he2e,
12'he67,
12'he83,
12'he7a,
12'he72,
12'he8b,
12'heae,
12'he9a,
12'he4b,
12'he10,
12'he0c,
12'he17,
12'he1f,
12'he2e,
12'he5b,
12'he9d,
12'hed4,
12'hf03,
12'hf23,
12'hf1f,
12'heff,
12'hebe,
12'he6c,
12'he2d,
12'he0c,
12'he0f,
12'he24,
12'he49,
12'hea9,
12'hf38,
12'hfb0,
12'hfd7,
12'hfb6,
12'hf75,
12'hf29,
12'heea,
12'hed6,
12'hee7,
12'hf0d,
12'hf28,
12'hf32,
12'hf72,
12'hfff,
12'h08b,
12'h0d1,
12'h0bc,
12'h076,
12'h02a,
12'hfeb,
12'hfe4,
12'h013,
12'h04d,
12'h072,
12'h06b,
12'h068,
12'h0b1,
12'h146,
12'h1e4,
12'h242,
12'h255,
12'h24f,
12'h248,
12'h22c,
12'h202,
12'h204,
12'h257,
12'h2b5,
12'h2dd,
12'h2eb,
12'h317,
12'h359,
12'h37f,
12'h362,
12'h308,
12'h2a8,
12'h25d,
12'h22d,
12'h225,
12'h236,
12'h24b,
12'h254,
12'h245,
12'h225,
12'h1fe,
12'h1d9,
12'h1bb,
12'h18f,
12'h158,
12'h125,
12'h0f2,
12'h0c6,
12'h0af,
12'h0aa,
12'h09d,
12'h073,
12'h03d,
12'h01d,
12'h013,
12'h00d,
12'hff8,
12'hfc1,
12'hf6b,
12'hef8,
12'he9a,
12'he8a,
12'heb4,
12'hef1,
12'hf18,
12'hf18,
12'hf0c,
12'hee9,
12'hecb,
12'hed6,
12'hefd,
12'hf0f,
12'hec6,
12'he53,
12'he12,
12'he11,
12'he3c,
12'he7c,
12'heb2,
12'heca,
12'hebd,
12'he94,
12'he84,
12'hebe,
12'hf1b,
12'hf49,
12'hf38,
12'hf0b,
12'hed4,
12'he9a,
12'he70,
12'he8c,
12'hef8,
12'hf60,
12'hf77,
12'hf55,
12'hf47,
12'hf6c,
12'hfae,
12'hfe6,
12'hff8,
12'hfdf,
12'hfaa,
12'hf67,
12'hf2b,
12'hf32,
12'hf98,
12'h027,
12'h08b,
12'h09b,
12'h078,
12'h056,
12'h03d,
12'h045,
12'h086,
12'h0f2,
12'h156,
12'h17d,
12'h164,
12'h132,
12'h114,
12'h112,
12'h10f,
12'h10f,
12'h126,
12'h143,
12'h137,
12'h0f5,
12'h0bc,
12'h0b5,
12'h0cf,
12'h0e1,
12'h0d4,
12'h0c3,
12'h0b8,
12'h0af,
12'h0a7,
12'h0af,
12'h0d6,
12'h105,
12'h106,
12'h0b5,
12'h03a,
12'hfd8,
12'hfac,
12'hfb2,
12'hfcc,
12'hff1,
12'h005,
12'hfe4,
12'hfac,
12'hf8f,
12'hf7e,
12'hf50,
12'hf02,
12'heb4,
12'he81,
12'he5f,
12'he46,
12'he48,
12'he6d,
12'he9e,
12'heb5,
12'hea3,
12'he83,
12'he75,
12'he76,
12'he6f,
12'he5c,
12'he50,
12'he64,
12'he90,
12'heb1,
12'hebe,
12'hec6,
12'hedb,
12'hefb,
12'hf1f,
12'hf2e,
12'hf10,
12'heea,
12'hec6,
12'he8a,
12'he44,
12'he13,
12'he15,
12'he42,
12'he9f,
12'hf23,
12'hf96,
12'hfdf,
12'hff1,
12'hfd7,
12'hfb4,
12'hf91,
12'hf64,
12'hf24,
12'hede,
12'heb2,
12'heb8,
12'hefe,
12'hf85,
12'h033,
12'h0d0,
12'h123,
12'h111,
12'h0c8,
12'h084,
12'h03b,
12'hfec,
12'hfaf,
12'hf97,
12'hfae,
12'hfe2,
12'h04d,
12'h106,
12'h1de,
12'h286,
12'h2ae,
12'h26f,
12'h236,
12'h222,
12'h203,
12'h1cb,
12'h1af,
12'h1d5,
12'h212,
12'h23c,
12'h26d,
12'h2d1,
12'h344,
12'h36b,
12'h336,
12'h2dc,
12'h287,
12'h22e,
12'h1f9,
12'h20e,
12'h230,
12'h224,
12'h1e8,
12'h1aa,
12'h192,
12'h180,
12'h164,
12'h153,
12'h159,
12'h15e,
12'h131,
12'h0de,
12'h0a7,
12'h093,
12'h06c,
12'h027,
12'hfea,
12'hfc7,
12'hfcb,
12'hfea,
12'h00b,
12'h011,
12'hfd2,
12'hf50,
12'heb2,
12'he3d,
12'he2a,
12'he5d,
12'heaa,
12'hefc,
12'hf3f,
12'hf68,
12'hf5d,
12'hf29,
12'hf0e,
12'hf12,
12'hefa,
12'he9a,
12'he20,
12'hde9,
12'he0b,
12'he57,
12'he9e,
12'hed4,
12'hef9,
12'hefc,
12'hecf,
12'he86,
12'he70,
12'heb1,
12'hf0a,
12'hf49,
12'hf5e,
12'hf48,
12'hf06,
12'heb7,
12'heaa,
12'hef2,
12'hf5d,
12'hf9f,
12'hf95,
12'hf78,
12'hf82,
12'hfb1,
12'hfe2,
12'hff4,
12'hfe0,
12'hfb8,
12'hf75,
12'hf25,
12'hf1c,
12'hf8b,
12'h034,
12'h0a2,
12'h0a9,
12'h085,
12'h076,
12'h079,
12'h07d,
12'h095,
12'h0de,
12'h137,
12'h161,
12'h150,
12'h125,
12'h10d,
12'h0fc,
12'h0e1,
12'h0dc,
12'h101,
12'h132,
12'h131,
12'h0ef,
12'h0a5,
12'h08d,
12'h09f,
12'h0bc,
12'h0d8,
12'h0df,
12'h0d2,
12'h0c7,
12'h0cf,
12'h0e5,
12'h0e8,
12'h0d5,
12'h0af,
12'h068,
12'h01d,
12'hff0,
12'hfe9,
12'hffa,
12'hff7,
12'hfd8,
12'hfbb,
12'hfa1,
12'hf7b,
12'hf63,
12'hf61,
12'hf5c,
12'hf3d,
12'hefc,
12'hec0,
12'he9f,
12'he7e,
12'he59,
12'he3d,
12'he4e,
12'he92,
12'hec6,
12'hec5,
12'hea3,
12'he90,
12'he85,
12'he4c,
12'he12,
12'he20,
12'he5f,
12'he92,
12'he9b,
12'heac,
12'hf02,
12'hf6f,
12'hfa6,
12'hf93,
12'hf55,
12'hf0e,
12'hebd,
12'he68,
12'he34,
12'he38,
12'he58,
12'he7c,
12'heac,
12'hf06,
12'hf86,
12'hfdc,
12'hfe0,
12'hfb1,
12'hf7b,
12'hf53,
12'hf24,
12'hf04,
12'hefc,
12'hefb,
12'hf08,
12'hf30,
12'hf90,
12'h01c,
12'h0a1,
12'h0e1,
12'h0c3,
12'h079,
12'h031,
12'h003,
12'hfe9,
12'hfe4,
12'hff3,
12'h00e,
12'h028,
12'h04b,
12'h0b9,
12'h16c,
12'h20d,
12'h256,
12'h23a,
12'h1f8,
12'h1da,
12'h1e4,
12'h1e1,
12'h1d5,
12'h200,
12'h263,
12'h2ba,
12'h2e5,
12'h314,
12'h36c,
12'h3a4,
12'h375,
12'h2fc,
12'h27f,
12'h21f,
12'h1ed,
12'h1ed,
12'h209,
12'h222,
12'h21a,
12'h1fd,
12'h1f3,
12'h1f8,
12'h1f7,
12'h1db,
12'h1b3,
12'h191,
12'h15a,
12'h117,
12'h0d8,
12'h0a3,
12'h07d,
12'h059,
12'h03b,
12'h030,
12'h047,
12'h06a,
12'h06c,
12'h044,
12'hff3,
12'hf91,
12'hf33,
12'hee6,
12'hec7,
12'hec8,
12'heca,
12'hec3,
12'hec7,
12'hee0,
12'hefa,
12'hf07,
12'hf14,
12'hf27,
12'hf25,
12'hee8,
12'he81,
12'he38,
12'he2e,
12'he58,
12'he7e,
12'he89,
12'he91,
12'he93,
12'he8e,
12'he85,
12'hea2,
12'hee6,
12'hf19,
12'hf1d,
12'hef7,
12'hece,
12'hec1,
12'hece,
12'hef5,
12'hf33,
12'hf5e,
12'hf52,
12'hf27,
12'hf15,
12'hf45,
12'hf9a,
12'hfd9,
12'hfdb,
12'hfb6,
12'hfa3,
12'hf9f,
12'hf93,
12'hf91,
12'hfc4,
12'h01a,
12'h049,
12'h045,
12'h04a,
12'h076,
12'h0a4,
12'h0ac,
12'h0a1,
12'h0b3,
12'h0f2,
12'h123,
12'h119,
12'h0f4,
12'h0e3,
12'h0de,
12'h0d2,
12'h0d6,
12'h105,
12'h152,
12'h16b,
12'h129,
12'h0d3,
12'h09a,
12'h087,
12'h08e,
12'h09c,
12'h0a9,
12'h0a6,
12'h09d,
12'h0a2,
12'h0bf,
12'h0ee,
12'h104,
12'h0e2,
12'h095,
12'h036,
12'hfe5,
12'hfc3,
12'hfcd,
12'hff3,
12'h013,
12'h00c,
12'hfe1,
12'hf99,
12'hf55,
12'hf3c,
12'hf33,
12'hf1c,
12'hef7,
12'hecf,
12'heba,
12'heaa,
12'he94,
12'he7e,
12'he85,
12'heb2,
12'hec7,
12'he9c,
12'he67,
12'he69,
12'he96,
12'hec0,
12'heb5,
12'he93,
12'he90,
12'he91,
12'he86,
12'he83,
12'heb4,
12'hf19,
12'hf5e,
12'hf5b,
12'hf20,
12'hee7,
12'hec5,
12'he9f,
12'he69,
12'he2d,
12'he05,
12'hdfd,
12'he2e,
12'heaa,
12'hf49,
12'hfc9,
12'hff5,
12'hfd7,
12'hf95,
12'hf5a,
12'hf33,
12'hf09,
12'hede,
12'hebb,
12'heab,
12'hecc,
12'hf20,
12'hf90,
12'h003,
12'h059,
12'h07e,
12'h075,
12'h054,
12'h02d,
12'hff5,
12'hfb4,
12'hf9c,
12'hfc1,
12'h006,
12'h05f,
12'h0cd,
12'h14a,
12'h1bf,
12'h200,
12'h203,
12'h1fb,
12'h217,
12'h23e,
12'h234,
12'h203,
12'h1ee,
12'h21b,
12'h270,
12'h2b6,
12'h2e6,
12'h328,
12'h362,
12'h364,
12'h32b,
12'h2e3,
12'h299,
12'h24b,
12'h224,
12'h220,
12'h21d,
12'h204,
12'h1d8,
12'h1c1,
12'h1b7,
12'h19b,
12'h177,
12'h161,
12'h166,
12'h163,
12'h131,
12'h0e1,
12'h08e,
12'h04f,
12'h024,
12'h008,
12'hff4,
12'hfdc,
12'hfd5,
12'hfd7,
12'hfc9,
12'hfa2,
12'hf5d,
12'hef9,
12'he91,
12'he4a,
12'he2d,
12'he34,
12'he5f,
12'heb5,
12'hf1b,
12'hf5c,
12'hf48,
12'hf11,
12'hef4,
12'hee5,
12'hec4,
12'he75,
12'he3f,
12'he5d,
12'hea7,
12'hed5,
12'heda,
12'hee6,
12'heef,
12'hee3,
12'heba,
12'he9d,
12'hebc,
12'hf0b,
12'hf5b,
12'hf95,
12'hfba,
12'hfbb,
12'hf94,
12'hf58,
12'hf39,
12'hf56,
12'hf96,
12'hfd9,
12'h012,
12'h044,
12'h05a,
12'h054,
12'h03c,
12'h029,
12'h035,
12'h040,
12'h01d,
12'hfe4,
12'hfd2,
12'h012,
12'h07e,
12'h0d8,
12'h11b,
12'h144,
12'h14d,
12'h10d,
12'h0a6,
12'h087,
12'h0d6,
12'h15a,
12'h1ab,
12'h1a2,
12'h15e,
12'h10f,
12'h0d8,
12'h0cc,
12'h0f3,
12'h12f,
12'h14d,
12'h12f,
12'h0e8,
12'h0a4,
12'h087,
12'h08c,
12'h0a2,
12'h0b7,
12'h0a1,
12'h056,
12'h010,
12'hffd,
12'h007,
12'h00f,
12'h007,
12'hff7,
12'hfd1,
12'hf98,
12'hf5c,
12'hf26,
12'hf0b,
12'hf04,
12'hf0a,
12'hf16,
12'hf07,
12'hed1,
12'he9f,
12'he87,
12'he7a,
12'he6a,
12'he3f,
12'he0f,
12'hde0,
12'hda7,
12'hd83,
12'hd99,
12'hde8,
12'he32,
12'he4d,
12'he34,
12'he0d,
12'hdef,
12'hdcd,
12'hdac,
12'hd9b,
12'hda2,
12'hdb1,
12'hdca,
12'hdff,
12'he49,
12'he89,
12'hea1,
12'he99,
12'he94,
12'he99,
12'he9a,
12'he97,
12'he95,
12'hea6,
12'hed3,
12'hf11,
12'hf55,
12'hfa1,
12'hfeb,
12'h00f,
12'h00c,
12'hfff,
12'h002,
12'h01e,
12'h03e,
12'h05c,
12'h073,
12'h091,
12'h0bc,
12'h0e7,
12'h112,
12'h13b,
12'h15b,
12'h16c,
12'h171,
12'h188,
12'h1bf,
12'h1ff,
12'h223,
12'h21e,
12'h210,
12'h20b,
12'h20f,
12'h220,
12'h246,
12'h27e,
12'h2ac,
12'h2c0,
12'h2c0,
12'h2b2,
12'h29f,
12'h28a,
12'h26d,
12'h244,
12'h21a,
12'h203,
12'h203,
12'h20a,
12'h20b,
12'h20c,
12'h216,
12'h212,
12'h1ff,
12'h1ea,
12'h1d0,
12'h1b1,
12'h18b,
12'h168,
12'h14e,
12'h146,
12'h147,
12'h12f,
12'h103,
12'h0cf,
12'h0a3,
12'h082,
12'h070,
12'h072,
12'h07c,
12'h079,
12'h056,
12'h023,
12'hff5,
12'hfce,
12'hfa1,
12'hf76,
12'hf5c,
12'hf44,
12'hf32,
12'hf2a,
12'hf39,
12'hf51,
12'hf59,
12'hf51,
12'hf37,
12'hf08,
12'hec8,
12'he91,
12'he6b,
12'he5b,
12'he63,
12'he7a,
12'he98,
12'head,
12'heaf,
12'he97,
12'he76,
12'he5f,
12'he60,
12'he66,
12'he6b,
12'he77,
12'he84,
12'he8f,
12'he8a,
12'he90,
12'heb1,
12'hed8,
12'heea,
12'hee4,
12'hee1,
12'hee2,
12'hee1,
12'hecc,
12'hebd,
12'heca,
12'hee3,
12'hefd,
12'hf18,
12'hf45,
12'hf67,
12'hf70,
12'hf67,
12'hf61,
12'hf69,
12'hf75,
12'hf79,
12'hf73,
12'hf84,
12'hfa7,
12'hfd4,
12'h001,
12'h026,
12'h03c,
12'h02d,
12'h009,
12'hfe4,
12'hfd8,
12'hfec,
12'h010,
12'h02e,
12'h02a,
12'h01f,
12'h01a,
12'h01b,
12'h01e,
12'h01d,
12'h01b,
12'h014,
12'h006,
12'hff4,
12'hfe8,
12'hfe8,
12'hfe5,
12'hfd2,
12'hfb6,
12'hfa4,
12'hfab,
12'hfc3,
12'hfdb,
12'hff2,
12'hffc,
12'hffb,
12'hff4,
12'hfed,
12'hfee,
12'hff9,
12'h000,
12'hff9,
12'hff3,
12'hff6,
12'h001,
12'h010,
12'h016,
12'h01c,
12'h029,
12'h03a,
12'h04c,
12'h069,
12'h086,
12'h096,
12'h098,
12'h08d,
12'h07d,
12'h073,
12'h07a,
12'h08b,
12'h0ac,
12'h0d7,
12'h0fe,
12'h11b,
12'h12c,
12'h136,
12'h13d,
12'h144,
12'h146,
12'h147,
12'h13d,
12'h12d,
12'h118,
12'h101,
12'h0fa,
12'h10b,
12'h126,
12'h134,
12'h130,
12'h118,
12'h107,
12'h101,
12'h103,
12'h10a,
12'h102,
12'h0f2,
12'h0d8,
12'h0bd,
12'h0a9,
12'h0a2,
12'h0ad,
12'h0b9,
12'h0b7,
12'h0a5,
12'h090,
12'h07e,
12'h071,
12'h061,
12'h046,
12'h02f,
12'h020,
12'h01b,
12'h026,
12'h036,
12'h03c,
12'h038,
12'h033,
12'h02d,
12'h023,
12'h01a,
12'h00e,
12'hfff,
12'hff2,
12'hfe1,
12'hfd0,
12'hfcc,
12'hfd3,
12'hfe0,
12'hfe5,
12'hfd8,
12'hfbf,
12'hfac,
12'hf9b,
12'hf82,
12'hf68,
12'hf55,
12'hf43,
12'hf2e,
12'hf18,
12'hf00,
12'hef0,
12'hede,
12'hecb,
12'heba,
12'hea4,
12'he92,
12'he81,
12'he75,
12'he71,
12'he77,
12'he8a,
12'he9b,
12'hea7,
12'heb7,
12'hec7,
12'hed1,
12'heda,
12'hee1,
12'heed,
12'hefd,
12'hefc,
12'hef4,
12'hef4,
12'hef0,
12'heeb,
12'hef1,
12'hf01,
12'hf1a,
12'hf32,
12'hf41,
12'hf4d,
12'hf54,
12'hf60,
12'hf72,
12'hf80,
12'hf85,
12'hf8b,
12'hf99,
12'hfa4,
12'hfab,
12'hfbb,
12'hfd1,
12'hfe4,
12'hfeb,
12'hfea,
12'hff0,
12'h001,
12'h01d,
12'h037,
12'h049,
12'h05c,
12'h06e,
12'h078,
12'h079,
12'h078,
12'h078,
12'h079,
12'h080,
12'h082,
12'h085,
12'h08f,
12'h0a5,
12'h0bf,
12'h0cd,
12'h0d5,
12'h0d7,
12'h0db,
12'h0dd,
12'h0e3,
12'h0f7,
12'h10d,
12'h121,
12'h12a,
12'h12d,
12'h12d,
12'h129,
12'h127,
12'h12e,
12'h131,
12'h127,
12'h118,
12'h10c,
12'h104,
12'h104,
12'h10d,
12'h10f,
12'h108,
12'h0fc,
12'h0e5,
12'h0d6,
12'h0d2,
12'h0cd,
12'h0c5,
12'h0b5,
12'h0a2,
12'h08a,
12'h070,
12'h062,
12'h062,
12'h063,
12'h05e,
12'h04e,
12'h03a,
12'h030,
12'h02a,
12'h029,
12'h02d,
12'h034,
12'h031,
12'h01e,
12'h004,
12'hfef,
12'hfde,
12'hfd2,
12'hfce,
12'hfc4,
12'hfae,
12'hf93,
12'hf76,
12'hf63,
12'hf53,
12'hf45,
12'hf43,
12'hf3f,
12'hf37,
12'hf30,
12'hf27,
12'hf23,
12'hf1e,
12'hf20,
12'hf1f,
12'hf0e,
12'hefa,
12'hef2,
12'hef7,
12'hefd,
12'hf08,
12'hf18,
12'hf22,
12'hf28,
12'hf26,
12'hf23,
12'hf27,
12'hf2b,
12'hf30,
12'hf2f,
12'hf2a,
12'hf26,
12'hf29,
12'hf33,
12'hf44,
12'hf58,
12'hf68,
12'hf73,
12'hf85,
12'hf97,
12'hfa8,
12'hfc1,
12'hfdc,
12'hff9,
12'h012,
12'h023,
12'h02d,
12'h02a,
12'h029,
12'h031,
12'h03d,
12'h049,
12'h04d,
12'h04c,
12'h04a,
12'h048,
12'h048,
12'h049,
12'h04e,
12'h059,
12'h060,
12'h058,
12'h049,
12'h044,
12'h04c,
12'h05c,
12'h06a,
12'h072,
12'h074,
12'h072,
12'h06c,
12'h06d,
12'h070,
12'h073,
12'h07b,
12'h083,
12'h089,
12'h088,
12'h087,
12'h082,
12'h079,
12'h078,
12'h075,
12'h06d,
12'h064,
12'h05b,
12'h05a,
12'h061,
12'h069,
12'h06d,
12'h068,
12'h063,
12'h05e,
12'h052,
12'h04c,
12'h04c,
12'h04e,
12'h04e,
12'h04d,
12'h049,
12'h043,
12'h044,
12'h046,
12'h045,
12'h040,
12'h033,
12'h02b,
12'h025,
12'h01e,
12'h01c,
12'h015,
12'h00d,
12'h007,
12'h001,
12'hfff,
12'hfff,
12'h000,
12'h007,
12'h00d,
12'h00f,
12'h00a,
12'h005,
12'h009,
12'h00c,
12'h014,
12'h015,
12'h00f,
12'h007,
12'hffb,
12'hff3,
12'hff5,
12'hffd,
12'h003,
12'h008,
12'h00d,
12'h00d,
12'h009,
12'h007,
12'h006,
12'h006,
12'h003,
12'hffe,
12'hff7,
12'hff1,
12'hfee,
12'hfeb,
12'hfe6,
12'hfe0,
12'hfdd,
12'hfdc,
12'hfd7,
12'hfd2,
12'hfce,
12'hfc7,
12'hfc4,
12'hfbd,
12'hfb3,
12'hfaa,
12'hfa0,
12'hf98,
12'hf8f,
12'hf87,
12'hf83,
12'hf83,
12'hf8a,
12'hf8a,
12'hf8a,
12'hf8b,
12'hf86,
12'hf7f,
12'hf77,
12'hf6f,
12'hf6b,
12'hf67,
12'hf62,
12'hf60,
12'hf5c,
12'hf5d,
12'hf5d,
12'hf5e,
12'hf60,
12'hf5c,
12'hf5b,
12'hf52,
12'hf4b,
12'hf48,
12'hf45,
12'hf50,
12'hf56,
12'hf5d,
12'hf6a,
12'hf73,
12'hf7f,
12'hf8b,
12'hf97,
12'hfa7,
12'hfb4,
12'hfbc,
12'hfc0,
12'hfc6,
12'hfcb,
12'hfcd,
12'hfd4,
12'hfd8,
12'hfe1,
12'hfea,
12'hfec,
12'hff5,
12'h000,
12'h00c,
12'h017,
12'h021,
12'h02c,
12'h036,
12'h046,
12'h051,
12'h059,
12'h061,
12'h064,
12'h06e,
12'h07a,
12'h084,
12'h08a,
12'h08d,
12'h096,
12'h0a0,
12'h0a8,
12'h0b0,
12'h0b8,
12'h0c0,
12'h0c8,
12'h0cc,
12'h0d1,
12'h0d7,
12'h0dc,
12'h0e2,
12'h0e4,
12'h0e0,
12'h0d8,
12'h0d1,
12'h0d1,
12'h0d2,
12'h0d2,
12'h0d3,
12'h0d1,
12'h0d2,
12'h0d4,
12'h0d4,
12'h0d0,
12'h0c9,
12'h0c0,
12'h0b7,
12'h0ad,
12'h0a3,
12'h09b,
12'h092,
12'h089,
12'h081,
12'h078,
12'h070,
12'h06c,
12'h067,
12'h05c,
12'h052,
12'h04a,
12'h03c,
12'h02d,
12'h020,
12'h014,
12'h00a,
12'h000,
12'hffe,
12'hff9,
12'hff3,
12'hfeb,
12'hfdf,
12'hfd6,
12'hfc6,
12'hfbc,
12'hfb6,
12'hfae,
12'hfa6,
12'hf98,
12'hf91,
12'hf8b,
12'hf86,
12'hf86,
12'hf87,
12'hf89,
12'hf80,
12'hf77,
12'hf78,
12'hf78,
12'hf71,
12'hf66,
12'hf5d,
12'hf56,
12'hf4c,
12'hf40,
12'hf3b,
12'hf3b,
12'hf3d,
12'hf3e,
12'hf3e,
12'hf40,
12'hf45,
12'hf4a,
12'hf4a,
12'hf4d,
12'hf4f,
12'hf4f,
12'hf52,
12'hf57,
12'hf5f,
12'hf65,
12'hf70,
12'hf7b,
12'hf83,
12'hf8f,
12'hf9a,
12'hfa3,
12'hfad,
12'hfb2,
12'hfb5,
12'hfbd,
12'hfc4,
12'hfc6,
12'hfcc,
12'hfd4,
12'hfdc,
12'hfe5,
12'hfec,
12'hff2,
12'hff5,
12'hff6,
12'hffd,
12'h004,
12'h011,
12'h01f,
12'h026,
12'h02c,
12'h02f,
12'h031,
12'h038,
12'h03a,
12'h03d,
12'h043,
12'h045,
12'h045,
12'h046,
12'h045,
12'h047,
12'h04c,
12'h04b,
12'h04a,
12'h04a,
12'h04a,
12'h046,
12'h045,
12'h048,
12'h046,
12'h044,
12'h03f,
12'h03d,
12'h041,
12'h045,
12'h049,
12'h04c,
12'h04a,
12'h049,
12'h048,
12'h04a,
12'h04f,
12'h04e,
12'h04b,
12'h04a,
12'h04c,
12'h050,
12'h051,
12'h054,
12'h058,
12'h05b,
12'h05c,
12'h05b,
12'h05c,
12'h058,
12'h04e,
12'h043,
12'h03f,
12'h03a,
12'h033,
12'h031,
12'h02f,
12'h031,
12'h02e,
12'h02e,
12'h033,
12'h036,
12'h03b,
12'h03c,
12'h039,
12'h039,
12'h038,
12'h035,
12'h036,
12'h036,
12'h02f,
12'h02a,
12'h028,
12'h027,
12'h024,
12'h01e,
12'h01f,
12'h023,
12'h026,
12'h028,
12'h02d,
12'h030,
12'h02b,
12'h029,
12'h025,
12'h021,
12'h01f,
12'h01a,
12'h017,
12'h014,
12'h00e,
12'h007,
12'h005,
12'h008,
12'h006,
12'h006,
12'h002,
12'hfff,
12'hffd,
12'hff5,
12'hff0,
12'hfec,
12'hfe7,
12'hfe2,
12'hfdb,
12'hfd3,
12'hfc9,
12'hfc3,
12'hfb8,
12'hfac,
12'hfa5,
12'hf9b,
12'hf97,
12'hf96,
12'hf97,
12'hf96,
12'hf91,
12'hf89,
12'hf80,
12'hf7f,
12'hf80,
12'hf7e,
12'hf7e,
12'hf7c,
12'hf7c,
12'hf7b,
12'hf7b,
12'hf7c,
12'hf7d,
12'hf7e,
12'hf7f,
12'hf7f,
12'hf80,
12'hf82,
12'hf83,
12'hf87,
12'hf8d,
12'hf91,
12'hf97,
12'hf9f,
12'hfa6,
12'hfa9,
12'hfaa,
12'hfae,
12'hfb2,
12'hfb6,
12'hfba,
12'hfbf,
12'hfc4,
12'hfc7,
12'hfcd,
12'hfd0,
12'hfd7,
12'hfe3,
12'hfec,
12'hfef,
12'hff3,
12'hff9,
12'hffe,
12'h005,
12'h00f,
12'h015,
12'h018,
12'h01a,
12'h022,
12'h028,
12'h02a,
12'h02f,
12'h036,
12'h03e,
12'h046,
12'h04e,
12'h056,
12'h05a,
12'h059,
12'h05d,
12'h063,
12'h066,
12'h06a,
12'h06c,
12'h072,
12'h074,
12'h072,
12'h075,
12'h075,
12'h077,
12'h079,
12'h077,
12'h079,
12'h07b,
12'h07c,
12'h07c,
12'h07f,
12'h081,
12'h07c,
12'h077,
12'h072,
12'h06c,
12'h06d,
12'h06a,
12'h064,
12'h062,
12'h05b,
12'h052,
12'h051,
12'h052,
12'h053,
12'h054,
12'h050,
12'h04e,
12'h04b,
12'h044,
12'h042,
12'h03c,
12'h038,
12'h034,
12'h02f,
12'h02f,
12'h02c,
12'h026,
12'h022,
12'h01e,
12'h01d,
12'h01a,
12'h018,
12'h016,
12'h00f,
12'h00a,
12'h002,
12'hffb,
12'hff9,
12'hff6,
12'hff1,
12'hfec,
12'hfe6,
12'hfe1,
12'hfdc,
12'hfd8,
12'hfd3,
12'hfd1,
12'hfce,
12'hfc9,
12'hfc6,
12'hfbe,
12'hfbb,
12'hfb6,
12'hfae,
12'hfae,
12'hfae,
12'hfac,
12'hfac,
12'hfad,
12'hfab,
12'hfaa,
12'hfa6,
12'hfa2,
12'hfa2,
12'hf9f,
12'hf9d,
12'hf9a,
12'hf97,
12'hf9a,
12'hf9b,
12'hf9b,
12'hfa1,
12'hfaa,
12'hfae,
12'hfad,
12'hfaf,
12'hfaf,
12'hfaf,
12'hfb0,
12'hfaf,
12'hfb3,
12'hfb7,
12'hfb8,
12'hfb6,
12'hfbb,
12'hfbf,
12'hfc0,
12'hfc6,
12'hfc9,
12'hfce,
12'hfd3,
12'hfd6,
12'hfdc,
12'hfdb,
12'hfdc,
12'hfdf,
12'hfe4,
12'hfec,
12'hfee,
12'hfed,
12'hff1,
12'hff5,
12'hff4,
12'hff8,
12'hffe,
12'h000,
12'h001,
12'h001,
12'h004,
12'h009,
12'h00d,
12'h011,
12'h018,
12'h01c,
12'h01d,
12'h01f,
12'h023,
12'h027,
12'h02b,
12'h02e,
12'h02d,
12'h02d,
12'h02e,
12'h02e,
12'h033,
12'h037,
12'h034,
12'h02f,
12'h02d,
12'h02e,
12'h02f,
12'h02d,
12'h02f,
12'h031,
12'h02f,
12'h02f,
12'h02d,
12'h02d,
12'h02a,
12'h026,
12'h02b,
12'h02c,
12'h02b,
12'h02b,
12'h02b,
12'h02d,
12'h02c,
12'h02d,
12'h02e,
12'h031,
12'h033,
12'h033,
12'h033,
12'h032,
12'h032,
12'h033,
12'h033,
12'h033,
12'h034,
12'h02f,
12'h02b,
12'h02c,
12'h02c,
12'h02b,
12'h02a,
12'h02c,
12'h02b,
12'h02a,
12'h02b,
12'h02c,
12'h02d,
12'h02c,
12'h02c,
12'h02b,
12'h02a,
12'h02a,
12'h02a,
12'h02a,
12'h02a,
12'h027,
12'h022,
12'h021,
12'h022,
12'h021,
12'h01d,
12'h01a,
12'h01a,
12'h017,
12'h010,
12'h00b,
12'h009,
12'h004,
12'h000,
12'h000,
12'hffa,
12'hff7,
12'hff4,
12'hff1,
12'hff1,
12'hfee,
12'hfea,
12'hfea,
12'hfe9,
12'hfe0,
12'hfdb,
12'hfd7,
12'hfd2,
12'hfd1,
12'hfd0,
12'hfd0,
12'hfcd,
12'hfca,
12'hfc4,
12'hfc1,
12'hfbf,
12'hfb8,
12'hfb5,
12'hfb1,
12'hfad,
12'hfaa,
12'hfa6,
12'hfa6,
12'hfa8,
12'hfa3,
12'hfa2,
12'hfa6,
12'hfa6,
12'hfa4,
12'hfa0,
12'hfa0,
12'hfa1,
12'hfa0,
12'hfa3,
12'hfa7,
12'hfa9,
12'hfac,
12'hfab,
12'hfb1,
12'hfb5,
12'hfb4,
12'hfb5,
12'hfb6,
12'hfbd,
12'hfbf,
12'hfbe,
12'hfc6,
12'hfc9,
12'hfcd,
12'hfd1,
12'hfd4,
12'hfd8,
12'hfdb,
12'hfe0,
12'hfe3,
12'hfe9,
12'hfeb,
12'hfe9,
12'hfef,
12'hff7,
12'hffe,
12'h007,
12'h009,
12'h00f,
12'h014,
12'h017,
12'h01a,
12'h01d,
12'h022,
12'h026,
12'h02a,
12'h02d,
12'h031,
12'h034,
12'h033,
12'h038,
12'h03d,
12'h03e,
12'h03e,
12'h03f,
12'h03f,
12'h03e,
12'h044,
12'h048,
12'h048,
12'h048,
12'h048,
12'h049,
12'h048,
12'h049,
12'h049,
12'h048,
12'h048,
12'h047,
12'h04c,
12'h04f,
12'h04b,
12'h049,
12'h04a,
12'h04a,
12'h049,
12'h043,
12'h045,
12'h049,
12'h044,
12'h041,
12'h040,
12'h03f,
12'h03b,
12'h037,
12'h038,
12'h035,
12'h031,
12'h031,
12'h030,
12'h030,
12'h02e,
12'h027,
12'h023,
12'h024,
12'h024,
12'h020,
12'h01c,
12'h01b,
12'h017,
12'h012,
12'h012,
12'h012,
12'h00e,
12'h00a,
12'h006,
12'h001,
12'hffe,
12'hff8,
12'hff2,
12'hff1,
12'hfee,
12'hfe9,
12'hfe8,
12'hfe5,
12'hfe2,
12'hfe0,
12'hfda,
12'hfd9,
12'hfd9,
12'hfd8,
12'hfd7,
12'hfd7,
12'hfd3,
12'hfcf,
12'hfce,
12'hfcc,
12'hfcd,
12'hfcc,
12'hfcc,
12'hfcd,
12'hfcd,
12'hfcf,
12'hfce,
12'hfcf,
12'hfcf,
12'hfcd,
12'hfcc,
12'hfcc,
12'hfcb,
12'hfcc,
12'hfcb,
12'hfcc,
12'hfcc,
12'hfc9,
12'hfca,
12'hfca,
12'hfca,
12'hfcc,
12'hfcc,
12'hfcb,
12'hfcb,
12'hfcb,
12'hfcc,
12'hfd2,
12'hfd4,
12'hfd3,
12'hfd3,
12'hfd3,
12'hfd6,
12'hfd5,
12'hfd8,
12'hfde,
12'hfdf,
12'hfe0,
12'hfe4,
12'hfe7,
12'hfe8,
12'hfe7,
12'hfe7,
12'hfec,
12'hff3,
12'hff0,
12'hff4,
12'hffa,
12'hffb,
12'hffb,
12'hffb,
12'h000,
12'h001,
12'h001,
12'h007,
12'h00a,
12'h009,
12'h00a,
12'h009,
12'h00d,
12'h012,
12'h013,
12'h014,
12'h015,
12'h01a,
12'h01c,
12'h01b,
12'h01e,
12'h01d,
12'h01e,
12'h01e,
12'h01f,
12'h01e,
12'h01d,
12'h01d,
12'h01d,
12'h01d,
12'h01f,
12'h020,
12'h021,
12'h022,
12'h023,
12'h026,
12'h029,
12'h029,
12'h029,
12'h028,
12'h026,
12'h029,
12'h028,
12'h028,
12'h02a,
12'h02a,
12'h02a,
12'h028,
12'h02c,
12'h030,
12'h030,
12'h030,
12'h031,
12'h031,
12'h031,
12'h031,
12'h030,
12'h02f,
12'h02b,
12'h025,
12'h026,
12'h026,
12'h022,
12'h01c,
12'h01c,
12'h01e,
12'h01e,
12'h01d,
12'h01c,
12'h018,
12'h013,
12'h010,
12'h00d,
12'h00c,
12'h00b,
12'h009,
12'h005,
12'h003,
12'h003,
12'h002,
12'hfff,
12'hffa,
12'hffa,
12'hff9,
12'hffb,
12'hff8,
12'hff2,
12'hff1,
12'hff2,
12'hfef,
12'hfea,
12'hfe8,
12'hfe9,
12'hfe7,
12'hfe7,
12'hfe6,
12'hfe4,
12'hfe2,
12'hfdd,
12'hfde,
12'hfdd,
12'hfdd,
12'hfdc,
12'hfd6,
12'hfd5,
12'hfd5,
12'hfd5,
12'hfd5,
12'hfd5,
12'hfd6,
12'hfd5,
12'hfd4,
12'hfd3,
12'hfd3,
12'hfd3,
12'hfd4,
12'hfd4,
12'hfd3,
12'hfd4,
12'hfd5,
12'hfd5,
12'hfd4,
12'hfd4,
12'hfd4,
12'hfd4,
12'hfd7,
12'hfdc,
12'hfdd,
12'hfdd,
12'hfdd,
12'hfde,
12'hfdf,
12'hfe3,
12'hfe7,
12'hfe5,
12'hfe9,
12'hfef,
12'hff0,
12'hff0,
12'hff1,
12'hff6,
12'hff9,
12'hff9,
12'hfff,
12'h001,
12'h000,
12'h000,
12'h003,
12'h009,
12'h009,
12'h009,
12'h00a,
12'h00b,
12'h00b,
12'h00b,
12'h00c,
12'h011,
12'h016,
12'h014,
12'h015,
12'h016,
12'h015,
12'h015,
12'h016,
12'h018,
12'h017,
12'h015,
12'h015,
12'h019,
12'h01c,
12'h018,
12'h018,
12'h017,
12'h017,
12'h015,
12'h015,
12'h017,
12'h018,
12'h019,
12'h017,
12'h019,
12'h019,
12'h018,
12'h016,
12'h016,
12'h015,
12'h010,
12'h010,
12'h010,
12'h011,
12'h012,
12'h012,
12'h011,
12'h011,
12'h011,
12'h00f,
12'h010,
12'h010,
12'h00f,
12'h010,
12'h010,
12'h011,
12'h010,
12'h00e,
12'h00e,
12'h009,
12'h005,
12'h005,
12'h004,
12'h005,
12'h005,
12'h004,
12'h004,
12'h004,
12'h003,
12'hfff,
12'hffc,
12'h000,
12'hfff,
12'hffa,
12'hffe,
12'hfff,
12'hffb,
12'hffa,
12'hff9,
12'hffa,
12'hffa,
12'hff8,
12'hff7,
12'hff7,
12'hff2,
12'hfee,
12'hfef,
12'hff0,
12'hff0,
12'hff0,
12'hfef,
12'hfef,
12'hfed,
12'hfe7,
12'hfe4,
12'hfe5,
12'hfe5,
12'hfe4,
12'hfe5,
12'hfe3,
12'hfdd,
12'hfdd,
12'hfde,
12'hfde,
12'hfde,
12'hfde,
12'hfdf,
12'hfe0,
12'hfe0,
12'hfdf,
12'hfde,
12'hfdf,
12'hfe0,
12'hfdf,
12'hfdf,
12'hfe0,
12'hfe1,
12'hfe0,
12'hfe1,
12'hfe7,
12'hfea,
12'hfea,
12'hfea,
12'hfeb,
12'hfea,
12'hfe8,
12'hfeb,
12'hff1,
12'hff3,
12'hff5,
12'hff6,
12'hff6,
12'hff9,
12'hffd,
12'hffe,
12'h001,
12'h006,
12'h006,
12'h009,
12'h00e,
12'h00f,
12'h00e,
12'h00e,
12'h014,
12'h016,
12'h016,
12'h017,
12'h01b,
12'h01f,
12'h01f,
12'h01f,
12'h022,
12'h026,
12'h027,
12'h028,
12'h028,
12'h028,
12'h029,
12'h027,
12'h026,
12'h027,
12'h027,
12'h028,
12'h02c,
12'h02f,
12'h030,
12'h02f,
12'h02e,
12'h02e,
12'h02d,
12'h02e,
12'h02d,
12'h02d,
12'h02b,
12'h026,
12'h025,
12'h024,
12'h025,
12'h026,
12'h025,
12'h025,
12'h01f,
12'h01c,
12'h01c,
12'h01b,
12'h018,
12'h013,
12'h013,
12'h012,
12'h011,
12'h012,
12'h012,
12'h011,
12'h00c,
12'h008,
12'h008,
12'h005,
12'h001,
12'hfff,
12'hfff,
12'h000,
12'hfff,
12'hff8,
12'hff7,
12'hff8,
12'hff6,
12'hff2,
12'hfee,
12'hfed,
12'hfea,
12'hfe5,
12'hfe5,
12'hfe4,
12'hfdf,
12'hfde,
12'hfdd,
12'hfdc,
12'hfdb,
12'hfd7,
12'hfd4,
12'hfd5,
12'hfd5,
12'hfd5,
12'hfd5,
12'hfd4,
12'hfd5,
12'hfd6,
12'hfd6,
12'hfd6,
12'hfd6,
12'hfd7,
12'hfd7,
12'hfd5,
12'hfd5,
12'hfd6,
12'hfd7,
12'hfd7,
12'hfd9,
12'hfd9,
12'hfd7,
12'hfd7,
12'hfd8,
12'hfd8,
12'hfd9,
12'hfde,
12'hfe2,
12'hfe2,
12'hfe2,
12'hfe3,
12'hfe3,
12'hfe2,
12'hfe3,
12'hfe4,
12'hfe4,
12'hfe9,
12'hfec,
12'hfec,
12'hfed,
12'hfef,
12'hff5,
12'hff6,
12'hff8,
12'hffd,
12'h000,
12'h000,
12'h000,
12'h003,
12'h007,
12'h008,
12'h007,
12'h006,
12'h007,
12'h009,
12'h00f,
12'h012,
12'h013,
12'h018,
12'h01b,
12'h01a,
12'h019,
12'h01a,
12'h01f,
12'h022,
12'h022,
12'h021,
12'h021,
12'h022,
12'h022,
12'h028,
12'h02b,
12'h02a,
12'h02a,
12'h02a,
12'h029,
12'h028,
12'h027,
12'h026,
12'h027,
12'h027,
12'h026,
12'h026,
12'h026,
12'h026,
12'h026,
12'h026,
12'h021,
12'h01e,
12'h01e,
12'h01d,
12'h01d,
12'h01e,
12'h01d,
12'h01d,
12'h01d,
12'h01d,
12'h01b,
12'h01b,
12'h01c,
12'h01c,
12'h01b,
12'h01d,
12'h01e,
12'h019,
12'h014,
12'h014,
12'h014,
12'h012,
12'h012,
12'h013,
12'h012,
12'h011,
12'h00d,
12'h00a,
12'h00b,
12'h00a,
12'h009,
12'h009,
12'h009,
12'h008,
12'h009,
12'h005,
12'h001,
12'h002,
12'h001,
12'h000,
12'h000,
12'h000,
12'hffe,
12'hffa,
12'hffa,
12'hff9,
12'hff8,
12'hff9,
12'hff8,
12'hff8,
12'hff9,
12'hff9,
12'hff4,
12'hfef,
12'hff1,
12'hff1,
12'hfef,
12'hfef,
12'hfef,
12'hff0,
12'hff1,
12'hfec,
12'hfe7,
12'hfe9,
12'hfe9,
12'hfe7,
12'hfe8,
12'hfe8,
12'hfe8,
12'hfe6,
12'hfe2,
12'hfe0,
12'hfe1,
12'hfe0,
12'hfe1,
12'hfe2,
12'hfde,
12'hfda,
12'hfd9,
12'hfda,
12'hfd9,
12'hfd9,
12'hfd9,
12'hfd9,
12'hfd9,
12'hfd4,
12'hfd2,
12'hfd3,
12'hfd2,
12'hfd2,
12'hfd2,
12'hfd3,
12'hfd3,
12'hfd2,
12'hfd2,
12'hfd2,
12'hfd3,
12'hfd4,
12'hfd4,
12'hfd5,
12'hfd5,
12'hfd5,
12'hfd5,
12'hfd7,
12'hfdc,
12'hfde,
12'hfdd,
12'hfde,
12'hfdf,
12'hfdf,
12'hfe4,
12'hfe8,
12'hfe7,
12'hfe6,
12'hfea,
12'hff0,
12'hff0,
12'hff0,
12'hff1,
12'hff1,
12'hff5,
12'hff8,
12'hff8,
12'hffd,
12'h000,
12'h000,
12'h000,
12'h002,
12'h008,
12'h009,
12'h009,
12'h00e,
12'h011,
12'h011,
12'h010,
12'h014,
12'h019,
12'h018,
12'h01b,
12'h01f,
12'h020,
12'h021,
12'h021,
12'h027,
12'h028,
12'h027,
12'h028,
12'h027,
12'h02c,
12'h02f,
12'h02f,
12'h030,
12'h02e,
12'h02e,
12'h02f,
12'h031,
12'h035,
12'h036,
12'h036,
12'h037,
12'h036,
12'h035,
12'h035,
12'h035,
12'h034,
12'h034,
12'h035,
12'h034,
12'h034,
12'h036,
12'h035,
12'h032,
12'h032,
12'h02e,
12'h02b,
12'h02b,
12'h02a,
12'h02a,
12'h029,
12'h028,
12'h028,
12'h023,
12'h020,
12'h021,
12'h021,
12'h01c,
12'h018,
12'h018,
12'h015,
12'h010,
12'h00f,
12'h00d,
12'h00c,
12'h007,
12'h005,
12'h005,
12'h000,
12'hffd,
12'hffd,
12'hffd,
12'hff9,
12'hff5,
12'hff6,
12'hff4,
12'hfed,
12'hfec,
12'hfed,
12'hfec,
12'hfe8,
12'hfe5,
12'hfe5,
12'hfe4,
12'hfe0,
12'hfdc,
12'hfdd,
12'hfdc,
12'hfdc,
12'hfdc,
12'hfd6,
12'hfd4,
12'hfd6,
12'hfd7,
12'hfd5,
12'hfd5,
12'hfd6,
12'hfd7,
12'hfd6,
12'hfd5,
12'hfd3,
12'hfcf,
12'hfce,
12'hfce,
12'hfcf,
12'hfd0,
12'hfcf,
12'hfd0,
12'hfd1,
12'hfd0,
12'hfd1,
12'hfd3,
12'hfd8,
12'hfdb,
12'hfda,
12'hfd9,
12'hfd9,
12'hfda,
12'hfda,
12'hfd9,
12'hfde,
12'hfe3,
12'hfe3,
12'hfe4,
12'hfe7,
12'hfeb,
12'hfed,
12'hfed,
12'hfee,
12'hfee,
12'hfed,
12'hff1,
12'hff6,
12'hff6,
12'hff7,
12'hff8,
12'hffa,
12'hffc,
12'hffd,
12'hfff,
12'h000,
12'h000,
12'h000,
12'h004,
12'h006,
12'h005,
12'h006,
12'h006,
12'h006,
12'h007,
12'h006,
12'h007,
12'h00d,
12'h00f,
12'h00e,
12'h00f,
12'h00e,
12'h00e,
12'h00e,
12'h00d,
12'h00c,
12'h00d,
12'h00e,
12'h00e,
12'h010,
12'h013,
12'h015,
12'h016,
12'h016,
12'h015,
12'h014,
12'h014,
12'h015,
12'h015,
12'h014,
12'h015,
12'h015,
12'h015,
12'h013,
12'h013,
12'h014,
12'h014,
12'h012,
12'h012,
12'h013,
12'h013,
12'h012,
12'h012,
12'h012,
12'h013,
12'h013,
12'h011,
12'h011,
12'h010,
12'h011,
12'h012,
12'h015,
12'h019,
12'h01a,
12'h019,
12'h019,
12'h019,
12'h01a,
12'h019,
12'h01a,
12'h019,
12'h01a,
12'h019,
12'h019,
12'h019,
12'h017,
12'h012,
12'h013,
12'h019,
12'h014,
12'h011,
12'h016,
12'h019,
12'h016,
12'h012,
12'h012,
12'h013,
12'h013,
12'h012,
12'h011,
12'h010,
12'h012,
12'h012,
12'h00c,
12'h009,
12'h00a,
12'h00b,
12'h009,
12'h00a,
12'h008,
12'h002,
12'h001,
12'h002,
12'h000,
12'h001,
12'h002,
12'hffe,
12'hff9,
12'hff8,
12'hffa,
12'hff7,
12'hff2,
12'hff1,
12'hff2,
12'hff0,
12'hfec,
12'hfe9,
12'hfea,
12'hfea,
12'hfe7,
12'hfe2,
12'hfe1,
12'hfe2,
12'hfe2,
12'hfe1,
12'hfe0,
12'hfdd,
12'hfda,
12'hfda,
12'hfd9,
12'hfd9,
12'hfd7,
12'hfd8,
12'hfd6,
12'hfd2,
12'hfd2,
12'hfd2,
12'hfd1,
12'hfd2,
12'hfd3,
12'hfd1,
12'hfd2,
12'hfd2,
12'hfd3,
12'hfd4,
12'hfd3,
12'hfd2,
12'hfd5,
12'hfd9,
12'hfd9,
12'hfda,
12'hfdc,
12'hfdd,
12'hfdd,
12'hfdd,
12'hfdd,
12'hfdd,
12'hfdf,
12'hfe3,
12'hfe5,
12'hfe5,
12'hfe6,
12'hfe7,
12'hfeb,
12'hfed,
12'hfed,
12'hfee,
12'hfee,
12'hff1,
12'hff5,
12'hff5,
12'hff4,
12'hff9,
12'hfff,
12'hfff,
12'hffe,
12'h000,
12'h003,
12'h006,
12'h005,
12'h005,
12'h009,
12'h00d,
12'h00c,
12'h00d,
12'h00d,
12'h00e,
12'h014,
12'h014,
12'h014,
12'h014,
12'h016,
12'h015,
12'h018,
12'h01c,
12'h01d,
12'h01c,
12'h01c,
12'h01c,
12'h01c,
12'h01c,
12'h01d,
12'h021,
12'h024,
12'h025,
12'h025,
12'h024,
12'h023,
12'h024,
12'h023,
12'h023,
12'h024,
12'h022,
12'h022,
12'h023,
12'h023,
12'h021,
12'h021,
12'h021,
12'h021,
12'h01d,
12'h018,
12'h019,
12'h019,
12'h018,
12'h019,
12'h019,
12'h018,
12'h017,
12'h018,
12'h017,
12'h014,
12'h011,
12'h010,
12'h010,
12'h010,
12'h00f,
12'h00f,
12'h010,
12'h00f,
12'h00b,
12'h008,
12'h009,
12'h008,
12'h009,
12'h008,
12'h008,
12'h006,
12'h001,
12'h000,
12'h002,
12'h001,
12'h000,
12'h000,
12'hffe,
12'hff9,
12'hffa,
12'hffa,
12'hff9,
12'hff9,
12'hffa,
12'hff9,
12'hff9,
12'hffa,
12'hff5,
12'hff3,
12'hff7,
12'hff5,
12'hff2,
12'hff2,
12'hff2,
12'hff3,
12'hff2,
12'hff2,
12'hff3,
12'hff4,
12'hff4,
12'hff2,
12'hff3,
12'hff4,
12'hff4,
12'hff2,
12'hff2,
12'hff2,
12'hff3,
12'hff3,
12'hff3,
12'hff3,
12'hff4,
12'hff4,
12'hff4,
12'hff4,
12'hff4,
12'hff3,
12'hff4,
12'hff4,
12'hff4,
12'hff4,
12'hff5,
12'hff4,
12'hff4,
12'hff4,
12'hff4,
12'hff4,
12'hff4,
12'hff7,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffa,
12'hffa,
12'hffc,
12'hffb,
12'hffa,
12'hffb,
12'hffb,
12'hffa,
12'hffa,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffb,
12'hffc,
12'hffb,
12'hffa,
12'hffa,
12'hffa,
12'hffc,
12'h000,
12'h003,
12'h002,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h001,
12'h003,
12'h009,
12'h00b,
12'h00a,
12'h009,
12'h009,
12'h00a,
12'h00b,
12'h00b,
12'h00a,
12'h00a,
12'h00a,
12'h009,
12'h009,
12'h00a,
12'h00b,
12'h00a,
12'h00b,
12'h00f,
12'h012,
12'h012,
12'h014,
12'h015,
12'h014,
12'h014,
12'h014,
12'h013,
12'h011,
12'h011,
12'h012,
12'h013,
12'h013,
12'h00f,
12'h010,
12'h013,
12'h00f,
12'h00b,
12'h00c,
12'h00c,
12'h00b,
12'h00b,
12'h00b,
12'h00c,
12'h00b,
12'h00b,
12'h00c,
12'h00b,
12'h007,
12'h003,
12'h004,
12'h004,
12'h002,
12'h003,
12'h003,
12'h002,
12'h002,
12'h000,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hff6,
12'hff3,
12'hff4,
12'hff3,
12'hff4,
12'hff5,
12'hff4,
12'hff4,
12'hff4,
12'hff4,
12'hff3,
12'hff2,
12'hff3,
12'hff2,
12'hff2,
12'hff3,
12'hff2,
12'hff2,
12'hff2,
12'hff2,
12'hfef,
12'hfea,
12'hfea,
12'hfeb,
12'hfec,
12'hff1,
12'hff4,
12'hff4,
12'hff3,
12'hff3,
12'hff3,
12'hff3,
12'hff3,
12'hff3,
12'hff2,
12'hff3,
12'hff3,
12'hff3,
12'hff3,
12'hff3,
12'hff4,
12'hff3,
12'hff5,
12'hffa,
12'hffb,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffb,
12'hffc,
12'hffc,
12'hfff,
12'h002,
12'h002,
12'h002,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h001,
12'h002,
12'h003,
12'h003,
12'h006,
12'h00b,
12'h00b,
12'h00a,
12'h00a,
12'h00a,
12'h00a,
12'h00a,
12'h009,
12'h00a,
12'h00b,
12'h00b,
12'h00b,
12'h00b,
12'h00a,
12'h00a,
12'h00b,
12'h00b,
12'h00a,
12'h00b,
12'h00a,
12'h005,
12'h003,
12'h004,
12'h004,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h003,
12'h002,
12'h002,
12'h000,
12'hffb,
12'hffc,
12'hffc,
12'hffb,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffb,
12'hffa,
12'hffa,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffa,
12'hffa,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffa,
12'hffa,
12'hffa,
12'hffb,
12'hffc,
12'hffc,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffe,
12'h002,
12'h002,
12'h002,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h006,
12'h00a,
12'h00b,
12'h00b,
12'h00a,
12'h00b,
12'h00c,
12'h00b,
12'h00b,
12'h00a,
12'h00a,
12'h00a,
12'h009,
12'h00a,
12'h00a,
12'h00a,
12'h00a,
12'h00b,
12'h00b,
12'h00a,
12'h009,
12'h00b,
12'h00b,
12'h00b,
12'h00b,
12'h00b,
12'h00b,
12'h00a,
12'h00b,
12'h00b,
12'h00a,
12'h00b,
12'h00b,
12'h00b,
12'h00b,
12'h006,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h001,
12'h002,
12'h000,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffb,
12'hff9,
12'hff5,
12'hff7,
12'hff6,
12'hff3,
12'hff4,
12'hff3,
12'hff3,
12'hff4,
12'hff3,
12'hff3,
12'hff2,
12'hff2,
12'hff2,
12'hff4,
12'hff9,
12'hffc,
12'hffb,
12'hffb,
12'hffa,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffb,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffe,
12'h002,
12'h001,
12'h001,
12'h002,
12'h002,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h001,
12'h001,
12'h002,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h001,
12'hffd,
12'hffb,
12'hffc,
12'hffb,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffa,
12'hffa,
12'hffa,
12'hffb,
12'hffb,
12'hffb,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffa,
12'hff9,
12'hffa,
12'hffa,
12'hffa,
12'hffb,
12'hffa,
12'hffa,
12'h000,
12'h002,
12'h001,
12'h002,
12'h001,
12'h001,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h000,
12'h001,
12'h002,
12'h001,
12'h002,
12'h002,
12'h002,
12'h004,
12'h007,
12'h009,
12'h009,
12'h00a,
12'h009,
12'h009,
12'h00a,
12'h00a,
12'h00b,
12'h00b,
12'h00a,
12'h00b,
12'h00b,
12'h00a,
12'h00b,
12'h00b,
12'h00c,
12'h00c,
12'h00b,
12'h00c,
12'h00b,
12'h00b,
12'h00c,
12'h00c,
12'h00b,
12'h00b,
12'h00b,
12'h00b,
12'h00a,
12'h00b,
12'h00c,
12'h00b,
12'h00a,
12'h009,
12'h00b,
12'h009,
12'h004,
12'h002,
12'h002,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h000,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffb,
12'hffb,
12'hffc,
12'hff7,
12'hff3,
12'hff4,
12'hff3,
12'hff3,
12'hff2,
12'hff2,
12'hff1,
12'hfed,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfeb,
12'hfec,
12'hfee,
12'hfed,
12'hfed,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfed,
12'hfec,
12'hfec,
12'hfed,
12'hfed,
12'hfec,
12'hfec,
12'hfeb,
12'hfec,
12'hfed,
12'hfee,
12'hfef,
12'hff1,
12'hff6,
12'hff5,
12'hff4,
12'hff4,
12'hff4,
12'hff4,
12'hff4,
12'hff9,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hfff,
12'hffd,
12'hfff,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h005,
12'h005,
12'h005,
12'h008,
12'h00c,
12'h00b,
12'h00b,
12'h00b,
12'h00c,
12'h00c,
12'h00c,
12'h00c,
12'h00b,
12'h011,
12'h014,
12'h013,
12'h014,
12'h014,
12'h014,
12'h014,
12'h013,
12'h013,
12'h013,
12'h014,
12'h013,
12'h013,
12'h014,
12'h013,
12'h013,
12'h013,
12'h013,
12'h013,
12'h013,
12'h014,
12'h014,
12'h014,
12'h013,
12'h013,
12'h013,
12'h012,
12'h012,
12'h010,
12'h00b,
12'h00b,
12'h00b,
12'h00b,
12'h00b,
12'h00a,
12'h00b,
12'h00a,
12'h00b,
12'h00a,
12'h009,
12'h009,
12'h009,
12'h00a,
12'h008,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'hfff,
12'hffc,
12'hffc,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffc,
12'hffd,
12'hffb,
12'hffa,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hff9,
12'hff4,
12'hff3,
12'hff4,
12'hff3,
12'hff3,
12'hff2,
12'hff6,
12'hff9,
12'hff5,
12'hff2,
12'hff3,
12'hff3,
12'hff3,
12'hff3,
12'hff2,
12'hff2,
12'hff2,
12'hff3,
12'hff3,
12'hff3,
12'hff3,
12'hff2,
12'hff2,
12'hff2,
12'hff3,
12'hff4,
12'hff3,
12'hff4,
12'hff4,
12'hff5,
12'hff5,
12'hff5,
12'hff5,
12'hff5,
12'hff4,
12'hff4,
12'hff4,
12'hff4,
12'hff4,
12'hff5,
12'hff5,
12'hff5,
12'hff9,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hfff,
12'h001,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h003,
12'h004,
12'h004,
12'h005,
12'h00a,
12'h00b,
12'h00b,
12'h00c,
12'h00c,
12'h00b,
12'h00a,
12'h00a,
12'h009,
12'h009,
12'h00a,
12'h00a,
12'h009,
12'h00c,
12'h012,
12'h013,
12'h013,
12'h013,
12'h012,
12'h013,
12'h013,
12'h012,
12'h013,
12'h013,
12'h013,
12'h012,
12'h012,
12'h011,
12'h011,
12'h011,
12'h012,
12'h011,
12'h00e,
12'h00a,
12'h00a,
12'h009,
12'h009,
12'h009,
12'h008,
12'h009,
12'h009,
12'h00a,
12'h00a,
12'h00a,
12'h00a,
12'h005,
12'h002,
12'h002,
12'h002,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'hffc,
12'hff9,
12'hffb,
12'hffb,
12'hffa,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hff9,
12'hff4,
12'hff2,
12'hff2,
12'hff1,
12'hff1,
12'hff1,
12'hff2,
12'hff2,
12'hfef,
12'hfeb,
12'hfeb,
12'hfeb,
12'hfec,
12'hfec,
12'hfeb,
12'hfeb,
12'hfeb,
12'hfeb,
12'hfec,
12'hfec,
12'hfec,
12'hfed,
12'hfed,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfec,
12'hfeb,
12'hfeb,
12'hfeb,
12'hfeb,
12'hfeb,
12'hfed,
12'hff1,
12'hff3,
12'hff4,
12'hff5,
12'hff5,
12'hff6,
12'hff6,
12'hff5,
12'hff4,
12'hff6,
12'hff6,
12'hff8,
12'hffc,
12'hffd,
12'hffc,
12'hffd,
12'hffe,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hfff,
12'h002,
12'h003,
12'h003,
12'h004,
12'h005,
12'h004,
12'h004,
12'h005,
12'h004,
12'h007,
12'h00a,
12'h00b,
12'h00b,
12'h00a,
12'h009,
12'h00a,
12'h00a,
12'h00a,
12'h00a,
12'h00a,
12'h00b,
12'h00c,
12'h00d,
12'h00d,
12'h00c,
12'h00d,
12'h00d,
12'h00c,
12'h00c,
12'h00c,
12'h00d,
12'h00d,
12'h00c,
12'h00b,
12'h00c,
12'h00b,
12'h00a,
12'h00a,
12'h009,
12'h009,
12'h00b,
12'h00a,
12'h00a,
12'h00a,
12'h009,
12'h009,
12'h00a,
12'h00a,
12'h00a,
12'h00c,
12'h00d,
12'h00c,
12'h00c,
12'h00d,
12'h00c,
12'h00c,
12'h00b,
12'h00a,
12'h006,
12'h004,
12'h004,
12'h002,
12'h002,
12'h002,
12'h002,
12'h001,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h002,
12'h002,
12'h001,
12'h002,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'hfff,
12'hffd,
12'hffb,
12'hffa,
12'hff9,
12'hff9,
12'hff9,
12'hffa,
12'hffc,
12'hffa,
12'hffa,
12'hffa,
12'hffa,
12'hffb,
12'hffa,
12'hff9,
12'hff9,
12'hff9,
12'hff9,
12'hffb,
12'hffa,
12'hff9,
12'hff9,
12'hff9,
12'hff9,
12'hff9,
12'hffa,
12'hffa,
12'hff9,
12'hffb,
12'hffb,
12'hffa,
12'hffa,
12'hffc,
12'hffc,
12'hffa,
12'hffc,
12'hffe,
12'hffc,
12'hffe,
12'hfff,
12'hffe,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffb,
12'hffb,
12'hffd,
12'hffe,
12'hfff,
12'hffe,
12'hffd,
12'hffd,
12'hffe,
12'hfff,
12'hfff,
12'hffe,
12'hfff,
12'hfff,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hffd,
12'hffd,
12'hffe,
12'hfff,
12'hfff,
12'hffe,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffe,
12'hffd,
12'hffd,
12'hffe,
12'hfff,
12'h000,
12'h002,
12'h003,
12'h003,
12'h004,
12'h005,
12'h004,
12'h004,
12'h004,
12'h003,
12'h002,
12'h003,
12'h004,
12'h005,
12'h005,
12'h006,
12'h005,
12'h004,
12'h004,
12'h004,
12'h005,
12'h006,
12'h005,
12'h004,
12'h004,
12'h004,
12'h004,
12'h005,
12'h006,
12'h009,
12'h00b,
12'h00b,
12'h00b,
12'h00b,
12'h00a,
12'h00b,
12'h00b,
12'h00b,
12'h00c,
12'h00c,
12'h00b,
12'h00b,
12'h00a,
12'h00b,
12'h00d,
12'h00d,
12'h00c,
12'h00b,
12'h00a,
12'h009,
12'h008,
12'h006,
12'h003,
12'h002,
12'h003,
12'h004,
12'h003,
12'h003,
12'h005,
12'h004,
12'h004,
12'h004,
12'h003,
12'h002,
12'h004,
12'h004,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h001,
12'h000,
12'hfff,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffe,
12'hffd,
12'hffc,
12'hffb,
12'hffa,
12'hffb,
12'hffc,
12'hffc,
12'hffb,
12'hffa,
12'hff9,
12'hffa,
12'hffa,
12'hffb,
12'hffb,
12'hff8,
12'hff5,
12'hff5,
12'hff6,
12'hff7,
12'hff8,
12'hff8,
12'hff7,
12'hff7,
12'hff6,
12'hff6,
12'hff7,
12'hff8,
12'hff9,
12'hffa,
12'hff9,
12'hffa,
12'hffd,
12'hfff,
12'hfff,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hfff,
12'hffe,
12'hfff,
12'h000,
12'hfff,
12'hffe,
12'hfff,
12'hffe,
12'hffd,
12'hffc,
12'hffa,
12'hffb,
12'hffd,
12'hfff,
12'h000,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffe,
12'h001,
12'h002,
12'h003,
12'h005,
12'h004,
12'h003,
12'h004,
12'h005,
12'h005,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h005,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h002,
12'h001,
12'h001,
12'h001,
12'h002,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h005,
12'h005,
12'h005,
12'h005,
12'h005,
12'h003,
12'h003,
12'h003,
12'h003,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'hffd,
12'hffb,
12'hffa,
12'hffa,
12'hffb,
12'hffc,
12'hffe,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffe,
12'hffe,
12'hffc,
12'hffb,
12'hffa,
12'hffb,
12'hffc,
12'hffc,
12'hffd,
12'hffe,
12'hffe,
12'hfff,
12'h000,
12'hfff,
12'h000,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'h000,
12'h001,
12'h000,
12'h000,
12'h001,
12'h002,
12'h004,
12'h005,
12'h005,
12'h004,
12'h003,
12'h002,
12'h001,
12'h002,
12'h003,
12'h004,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h005,
12'h004,
12'h003,
12'h004,
12'h004,
12'h004,
12'h005,
12'h006,
12'h005,
12'h005,
12'h004,
12'h003,
12'h004,
12'h003,
12'h003,
12'h002,
12'h001,
12'h002,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h001,
12'h002,
12'h003,
12'h002,
12'h001,
12'h001,
12'h001,
12'h002,
12'h002,
12'h002,
12'h002,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h002,
12'h002,
12'h001,
12'h002,
12'h001,
12'hfff,
12'hffd,
12'hffc,
12'hffb,
12'hffb,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffb,
12'hffa,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffc,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffa,
12'hffb,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hffd,
12'hffe,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffe,
12'hfff,
12'hfff,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hfff,
12'hffe,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hfff,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hffe,
12'hfff,
12'hfff,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'h000,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h004,
12'h005,
12'h005,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h005,
12'h005,
12'h005,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h001,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'hfff,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffb,
12'hffd,
12'hffc,
12'hffc,
12'hffb,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffb,
12'hffb,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffb,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffb,
12'hffc,
12'hffc,
12'hffd,
12'hffe,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hfff,
12'h003,
12'h005,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h003,
12'h003,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'hfff,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hffe,
12'hffd,
12'hfff,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h005,
12'h004,
12'h005,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h004,
12'h003,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h000,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'h000,
12'h003,
12'h002,
12'h003,
12'h003,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h004,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'hfff,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'h000,
12'h000,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'h000,
12'h003,
12'h004,
12'h003,
12'h004,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h004,
12'h005,
12'h004,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h005,
12'h004,
12'h005,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h000,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hffd,
12'hffe,
12'hffe,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'h003,
12'h001,
12'hffe,
12'h001,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h002,
12'h003,
12'h003,
12'h002,
12'hffe,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffc,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffd,
12'hffe,
12'hffe,
12'hffd,
12'h001,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h004,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h004,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h004,
12'h003,
12'hfff,
12'hffd,
12'hffe,
12'hffe,
12'hffd,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffe,
12'hffe,
12'hffe,
12'hffd,
12'hffe,
12'hffe,
12'hffe,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffd,
12'h000,
12'h004,
12'h000,
12'h000,
12'h003,
12'h003,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h004,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h004,
12'h004,
12'h003,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h004,
12'h004,
12'h004,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'hfff,
12'hffc,
12'hffc,
12'hffb,
12'hffc,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffd,
12'hffc,
12'hffc,
12'hffc,
12'hffc,
12'hffd,
12'hffc,
12'hffd,
12'hffd,
12'h000,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h002,
12'h003,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h003,
12'h003,
12'h003,
12'h003,
12'h003,
12'h002,
12'h003,
12'h003,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h001,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h001,
12'h002,
12'h002,
12'h001,
12'h001,
12'h002,
12'h002,
12'h002,
12'h002,
12'h001,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h001,
12'h001,
12'h002,
12'h002,
12'h002,
12'h002,
12'h002,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h002,
12'h002,
12'h001,
12'h001,
12'h001,
12'h002,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h002,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h002,
12'h002,
12'h001,
12'h002,
12'h002,
12'h001,
12'h002,
12'h002,
12'h002,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h002,
12'h001,
12'h001,
12'h001,
12'h002,
12'h002,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h001,
12'h000,
12'h000,
12'h001
};

endpackage
