package obj_pkg;

localparam int NUM_OBJ = 4;
localparam int MAX_SIZE_Y = 64;
localparam int MAX_SIZE_X = 16;

localparam int ObjSizeX [NUM_OBJ-1:0] = {16, 16, 16, 16};
localparam int ObjSizeY [NUM_OBJ-1:0] = {64, 64, 16, 16};

localparam logic [NUM_OBJ-1:0][MAX_SIZE_Y-1:0][MAX_SIZE_X-1:0] Obj = {
  // object 3
  {
    {16'b1111111100000000},
    {16'b1111111100000000},
    {16'b1111111100000000},
    {16'b1111111100000000},
    {16'b1111111110000000},
    {16'b1111111110000000},
    {16'b1111111110000000},
    {16'b1111111110000000},
    {16'b1111111111000000},
    {16'b1111111111000000},
    {16'b1111111111000000},
    {16'b1111111111000000},
    {16'b1111111111100000},
    {16'b1111111111100000},
    {16'b1111111111100000},
    {16'b1111111111100000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111110000},
    {16'b1111111111100000},
    {16'b1111111111100000},
    {16'b1111111111100000},
    {16'b1111111111100000},
    {16'b1111111111000000},
    {16'b1111111111000000},
    {16'b1111111111000000},
    {16'b1111111111000000},
    {16'b1111111110000000},
    {16'b1111111110000000},
    {16'b1111111110000000},
    {16'b1111111110000000},
    {16'b1111111100000000},
    {16'b1111111100000000},
    {16'b1111111100000000},
    {16'b1111111100000000}
  },
  // object 2:
  {
    {16'b0000000011111111},
    {16'b0000000011111111},
    {16'b0000000011111111},
    {16'b0000000011111111},
    {16'b0000000111111111},
    {16'b0000000111111111},
    {16'b0000000111111111},
    {16'b0000000111111111},
    {16'b0000001111111111},
    {16'b0000001111111111},
    {16'b0000001111111111},
    {16'b0000001111111111},
    {16'b0000011111111111},
    {16'b0000011111111111},
    {16'b0000011111111111},
    {16'b0000011111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000111111111111},
    {16'b0000011111111111},
    {16'b0000011111111111},
    {16'b0000011111111111},
    {16'b0000011111111111},
    {16'b0000001111111111},
    {16'b0000001111111111},
    {16'b0000001111111111},
    {16'b0000001111111111},
    {16'b0000000111111111},
    {16'b0000000111111111},
    {16'b0000000111111111},
    {16'b0000000111111111},
    {16'b0000000011111111},
    {16'b0000000011111111},
    {16'b0000000011111111},
    {16'b0000000011111111}
  },
  // object 1:
  {
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000011111100000},
    {16'b0001111111111000},
    {16'b0011111111111100},
    {16'b0111111111111110},
    {16'b0111111111111110},
    {16'b1111111111111111},
    {16'b1111111111111111},
    {16'b1111111111111111},
    {16'b1111111111111111},
    {16'b1111111111111111},
    {16'b1111111111111111},
    {16'b0111111111111110},
    {16'b0111111111111110},
    {16'b0011111111111100},
    {16'b0001111111111000},
    {16'b0000011111100000}
  },
  // object 0
  {
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000000000000000},
    {16'b0000011111100000},
    {16'b0001111111111000},
    {16'b0011111111111100},
    {16'b0111111111111110},
    {16'b0111111111111110},
    {16'b1111111111111111},
    {16'b1111111111111111},
    {16'b1111111001111111},
    {16'b1111111001111111},
    {16'b1111111111111111},
    {16'b1111111111111111},
    {16'b0111111111111110},
    {16'b0111111111111110},
    {16'b0011111111111100},
    {16'b0001111111111000},
    {16'b0000011111100000}
  }
  };


endpackage
